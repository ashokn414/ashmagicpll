* NGSPICE file created from mux.ext - technology: sky130A


* Top level circuit mux

X0 i1 se vdd vdd sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X1 out se i1 vdd sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X2 i2 se out gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 i1 se gnd gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 out i1 i1 gnd sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 i2 i1 out vdd sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
.end

