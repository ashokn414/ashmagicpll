magic
tech sky130A
timestamp 1605617331
<< psubdiff >>
rect 70 1382 140 1402
rect 70 1352 90 1382
rect 120 1352 140 1382
rect 70 1332 140 1352
rect 170 1382 240 1402
rect 170 1352 190 1382
rect 220 1352 240 1382
rect 170 1332 240 1352
rect 270 1382 340 1402
rect 270 1352 290 1382
rect 320 1352 340 1382
rect 270 1332 340 1352
rect 370 1382 440 1402
rect 370 1352 390 1382
rect 420 1352 440 1382
rect 370 1332 440 1352
rect 470 1382 540 1402
rect 470 1352 490 1382
rect 520 1352 540 1382
rect 470 1332 540 1352
rect 570 1382 640 1402
rect 570 1352 590 1382
rect 620 1352 640 1382
rect 570 1332 640 1352
rect 670 1382 740 1402
rect 670 1352 690 1382
rect 720 1352 740 1382
rect 670 1332 740 1352
rect 770 1382 848 1402
rect 770 1352 790 1382
rect 820 1352 848 1382
rect 770 1332 848 1352
rect 878 1382 958 1402
rect 878 1352 898 1382
rect 928 1352 958 1382
rect 878 1332 958 1352
rect 988 1382 1071 1402
rect 988 1352 1021 1382
rect 1051 1352 1071 1382
rect 988 1332 1071 1352
rect 1101 1382 1191 1402
rect 1101 1352 1141 1382
rect 1171 1352 1191 1382
rect 1101 1332 1191 1352
rect 1221 1382 1291 1402
rect 1221 1352 1241 1382
rect 1271 1352 1291 1382
rect 1221 1332 1291 1352
rect 1321 1382 1395 1402
rect 1321 1352 1341 1382
rect 1371 1352 1395 1382
rect 1321 1332 1395 1352
rect 1425 1382 1495 1402
rect 1425 1352 1445 1382
rect 1475 1352 1495 1382
rect 1425 1332 1495 1352
rect 1553 1382 1623 1402
rect 1553 1352 1573 1382
rect 1603 1352 1623 1382
rect 1553 1332 1623 1352
rect 1653 1382 1723 1402
rect 1653 1352 1673 1382
rect 1703 1352 1723 1382
rect 1653 1332 1723 1352
rect 1753 1382 1823 1402
rect 1753 1352 1773 1382
rect 1803 1352 1823 1382
rect 1753 1332 1823 1352
rect 1853 1382 1923 1402
rect 1853 1352 1873 1382
rect 1903 1352 1923 1382
rect 1853 1332 1923 1352
rect 1953 1382 2023 1402
rect 1953 1352 1973 1382
rect 2003 1352 2023 1382
rect 1953 1332 2023 1352
rect 2053 1382 2123 1402
rect 2053 1352 2073 1382
rect 2103 1352 2123 1382
rect 2053 1332 2123 1352
rect 2153 1382 2223 1402
rect 2153 1352 2173 1382
rect 2203 1352 2223 1382
rect 2153 1332 2223 1352
rect 2253 1382 2331 1402
rect 2253 1352 2273 1382
rect 2303 1352 2331 1382
rect 2253 1332 2331 1352
rect 2361 1382 2441 1402
rect 2361 1352 2381 1382
rect 2411 1352 2441 1382
rect 2361 1332 2441 1352
rect 2471 1382 2554 1402
rect 2471 1352 2504 1382
rect 2534 1352 2554 1382
rect 2471 1332 2554 1352
rect 2584 1382 2674 1402
rect 2584 1352 2624 1382
rect 2654 1352 2674 1382
rect 2584 1332 2674 1352
rect 2704 1382 2774 1402
rect 2704 1352 2724 1382
rect 2754 1352 2774 1382
rect 2704 1332 2774 1352
rect 2804 1382 2878 1402
rect 2804 1352 2824 1382
rect 2854 1352 2878 1382
rect 2804 1332 2878 1352
rect 2908 1382 2978 1402
rect 2908 1352 2928 1382
rect 2958 1352 2978 1382
rect 2908 1332 2978 1352
rect 3039 1382 3109 1402
rect 3039 1352 3059 1382
rect 3089 1352 3109 1382
rect 3039 1332 3109 1352
rect 3139 1382 3209 1402
rect 3139 1352 3159 1382
rect 3189 1352 3209 1382
rect 3139 1332 3209 1352
rect 3239 1382 3309 1402
rect 3239 1352 3259 1382
rect 3289 1352 3309 1382
rect 3239 1332 3309 1352
rect 3339 1382 3409 1402
rect 3339 1352 3359 1382
rect 3389 1352 3409 1382
rect 3339 1332 3409 1352
rect 3439 1382 3509 1402
rect 3439 1352 3459 1382
rect 3489 1352 3509 1382
rect 3439 1332 3509 1352
rect 3539 1382 3609 1402
rect 3539 1352 3559 1382
rect 3589 1352 3609 1382
rect 3539 1332 3609 1352
rect 3639 1382 3709 1402
rect 3639 1352 3659 1382
rect 3689 1352 3709 1382
rect 3639 1332 3709 1352
rect 3739 1382 3817 1402
rect 3739 1352 3759 1382
rect 3789 1352 3817 1382
rect 3739 1332 3817 1352
rect 3847 1382 3927 1402
rect 3847 1352 3867 1382
rect 3897 1352 3927 1382
rect 3847 1332 3927 1352
rect 3957 1382 4040 1402
rect 3957 1352 3990 1382
rect 4020 1352 4040 1382
rect 3957 1332 4040 1352
rect 4070 1382 4160 1402
rect 4070 1352 4110 1382
rect 4140 1352 4160 1382
rect 4070 1332 4160 1352
rect 4190 1382 4260 1402
rect 4190 1352 4210 1382
rect 4240 1352 4260 1382
rect 4190 1332 4260 1352
rect 4290 1382 4364 1402
rect 4290 1352 4310 1382
rect 4340 1352 4364 1382
rect 4290 1332 4364 1352
rect 4394 1382 4464 1402
rect 4394 1352 4414 1382
rect 4444 1352 4464 1382
rect 4394 1332 4464 1352
<< psubdiffcont >>
rect 90 1352 120 1382
rect 190 1352 220 1382
rect 290 1352 320 1382
rect 390 1352 420 1382
rect 490 1352 520 1382
rect 590 1352 620 1382
rect 690 1352 720 1382
rect 790 1352 820 1382
rect 898 1352 928 1382
rect 1021 1352 1051 1382
rect 1141 1352 1171 1382
rect 1241 1352 1271 1382
rect 1341 1352 1371 1382
rect 1445 1352 1475 1382
rect 1573 1352 1603 1382
rect 1673 1352 1703 1382
rect 1773 1352 1803 1382
rect 1873 1352 1903 1382
rect 1973 1352 2003 1382
rect 2073 1352 2103 1382
rect 2173 1352 2203 1382
rect 2273 1352 2303 1382
rect 2381 1352 2411 1382
rect 2504 1352 2534 1382
rect 2624 1352 2654 1382
rect 2724 1352 2754 1382
rect 2824 1352 2854 1382
rect 2928 1352 2958 1382
rect 3059 1352 3089 1382
rect 3159 1352 3189 1382
rect 3259 1352 3289 1382
rect 3359 1352 3389 1382
rect 3459 1352 3489 1382
rect 3559 1352 3589 1382
rect 3659 1352 3689 1382
rect 3759 1352 3789 1382
rect 3867 1352 3897 1382
rect 3990 1352 4020 1382
rect 4110 1352 4140 1382
rect 4210 1352 4240 1382
rect 4310 1352 4340 1382
rect 4414 1352 4444 1382
<< locali >>
rect -111 1990 100 2020
rect -111 660 -61 1990
rect 2839 1510 2869 1681
rect 2839 1480 4630 1510
rect 0 1382 4504 1410
rect 0 1352 90 1382
rect 120 1352 190 1382
rect 220 1352 290 1382
rect 320 1352 390 1382
rect 420 1352 490 1382
rect 520 1352 590 1382
rect 620 1352 690 1382
rect 720 1352 790 1382
rect 820 1352 898 1382
rect 928 1352 1021 1382
rect 1051 1352 1141 1382
rect 1171 1352 1241 1382
rect 1271 1352 1341 1382
rect 1371 1352 1445 1382
rect 1475 1352 1573 1382
rect 1603 1352 1673 1382
rect 1703 1352 1773 1382
rect 1803 1352 1873 1382
rect 1903 1352 1973 1382
rect 2003 1352 2073 1382
rect 2103 1352 2173 1382
rect 2203 1352 2273 1382
rect 2303 1352 2381 1382
rect 2411 1352 2504 1382
rect 2534 1352 2624 1382
rect 2654 1352 2724 1382
rect 2754 1352 2824 1382
rect 2854 1352 2928 1382
rect 2958 1352 3059 1382
rect 3089 1352 3159 1382
rect 3189 1352 3259 1382
rect 3289 1352 3359 1382
rect 3389 1352 3459 1382
rect 3489 1352 3559 1382
rect 3589 1352 3659 1382
rect 3689 1352 3759 1382
rect 3789 1352 3867 1382
rect 3897 1352 3990 1382
rect 4020 1352 4110 1382
rect 4140 1352 4210 1382
rect 4240 1352 4310 1382
rect 4340 1352 4414 1382
rect 4444 1352 4504 1382
rect 0 1284 4504 1352
rect 1470 872 1510 880
rect 2980 875 3020 880
rect 4590 875 4630 1480
rect 1433 865 1510 872
rect 1433 843 1480 865
rect 1500 843 1510 865
rect 1433 840 1510 843
rect 2916 865 3020 875
rect 2916 843 2990 865
rect 3010 843 3020 865
rect 4402 844 4630 875
rect 2916 840 3020 843
rect 1470 830 1510 840
rect 2980 830 3020 840
rect -111 640 -100 660
rect -74 640 -61 660
rect -111 630 -61 640
<< viali >>
rect 1480 843 1500 865
rect 2990 843 3010 865
rect -100 640 -74 660
<< metal1 >>
rect 1470 865 1510 880
rect 1470 843 1480 865
rect 1500 843 1510 865
rect 1470 830 1510 843
rect 2980 865 3020 880
rect 2980 843 2990 865
rect 3010 843 3020 865
rect 2980 830 3020 843
rect -111 660 -61 670
rect -111 640 -100 660
rect -74 640 23 660
rect -111 630 23 640
rect 1480 630 1510 830
rect 2990 630 3020 830
use freq_div_2pll  freq_div_2pll_0 ~/Desktop/vsd/magic_exp/ashmagicpll
timestamp 1605609062
transform -1 0 1480 0 -1 300
box -65 -1034 1480 300
use freq_div_2pll  freq_div_2pll_1
timestamp 1605609062
transform -1 0 2963 0 -1 300
box -65 -1034 1480 300
use pfdpll  pfdpll_0 ~/Desktop/vsd/magic_exp/ashmagicpll
timestamp 1605604810
transform 1 0 130 0 1 4011
box -130 -2441 1390 610
use freq_div_2pll  freq_div_2pll_2
timestamp 1605609062
transform -1 0 4449 0 -1 300
box -65 -1034 1480 300
use vcopll  vcopll_0 ~/Desktop/vsd/magic_exp/ashmagicpll
timestamp 1605609241
transform 0 1 3109 -1 0 3131
box -20 -549 1500 90
<< labels >>
rlabel space 2847 1691 2863 1702 1 fvco_8
<< end >>
