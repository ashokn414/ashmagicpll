magic
tech sky130A
timestamp 1605510618
<< nwell >>
rect -10 -190 510 118
<< nmos >>
rect 90 -440 105 -398
rect 270 -440 285 -398
rect 360 -440 375 -398
<< pmos >>
rect 90 -144 105 -32
rect 270 -144 285 -32
rect 355 -144 370 -32
<< ndiff >>
rect 30 -408 90 -398
rect 30 -432 38 -408
rect 62 -432 90 -408
rect 30 -440 90 -432
rect 105 -406 270 -398
rect 105 -432 128 -406
rect 154 -432 208 -406
rect 234 -432 270 -406
rect 105 -440 270 -432
rect 285 -406 360 -398
rect 285 -432 308 -406
rect 334 -432 360 -406
rect 285 -440 360 -432
rect 375 -406 440 -398
rect 375 -432 408 -406
rect 434 -432 440 -406
rect 375 -440 440 -432
<< pdiff >>
rect 30 -80 90 -32
rect 30 -120 40 -80
rect 70 -120 90 -80
rect 30 -144 90 -120
rect 105 -80 160 -32
rect 105 -120 125 -80
rect 155 -120 160 -80
rect 105 -144 160 -120
rect 200 -80 270 -32
rect 200 -120 205 -80
rect 235 -120 270 -80
rect 200 -144 270 -120
rect 285 -80 355 -32
rect 285 -120 305 -80
rect 335 -120 355 -80
rect 285 -144 355 -120
rect 370 -80 440 -32
rect 370 -120 404 -80
rect 434 -120 440 -80
rect 370 -144 440 -120
<< ndiffc >>
rect 38 -432 62 -408
rect 128 -432 154 -406
rect 208 -432 234 -406
rect 308 -432 334 -406
rect 408 -432 434 -406
<< pdiffc >>
rect 40 -120 70 -80
rect 125 -120 155 -80
rect 205 -120 235 -80
rect 305 -120 335 -80
rect 404 -120 434 -80
<< psubdiff >>
rect 10 -510 490 -500
rect 10 -550 30 -510
rect 70 -550 110 -510
rect 150 -550 190 -510
rect 230 -550 270 -510
rect 310 -550 350 -510
rect 390 -550 430 -510
rect 470 -550 490 -510
rect 10 -560 490 -550
<< nsubdiff >>
rect 10 88 490 98
rect 10 48 30 88
rect 70 48 110 88
rect 150 48 190 88
rect 230 48 270 88
rect 310 48 350 88
rect 390 48 430 88
rect 470 48 490 88
rect 10 38 490 48
<< psubdiffcont >>
rect 30 -550 70 -510
rect 110 -550 150 -510
rect 190 -550 230 -510
rect 270 -550 310 -510
rect 350 -550 390 -510
rect 430 -550 470 -510
<< nsubdiffcont >>
rect 30 48 70 88
rect 110 48 150 88
rect 190 48 230 88
rect 270 48 310 88
rect 350 48 390 88
rect 430 48 470 88
<< poly >>
rect 90 -32 105 -12
rect 270 -32 285 -12
rect 355 -32 370 -12
rect 90 -180 105 -144
rect 270 -180 285 -144
rect 70 -193 110 -180
rect 70 -220 79 -193
rect 102 -220 110 -193
rect 70 -230 110 -220
rect 260 -194 300 -180
rect 260 -216 270 -194
rect 290 -216 300 -194
rect 260 -230 300 -216
rect 90 -313 105 -230
rect 355 -270 370 -144
rect 270 -285 370 -270
rect 270 -310 285 -285
rect 70 -324 110 -313
rect 70 -349 79 -324
rect 102 -349 110 -324
rect 70 -360 110 -349
rect 260 -321 300 -310
rect 260 -347 268 -321
rect 294 -347 300 -321
rect 260 -360 300 -347
rect 350 -324 390 -310
rect 350 -346 360 -324
rect 380 -346 390 -324
rect 350 -360 390 -346
rect 90 -398 105 -360
rect 270 -398 285 -360
rect 360 -398 375 -360
rect 90 -460 105 -440
rect 270 -460 285 -440
rect 360 -460 375 -440
<< polycont >>
rect 79 -220 102 -193
rect 270 -216 290 -194
rect 79 -349 102 -324
rect 268 -347 294 -321
rect 360 -346 380 -324
<< locali >>
rect 0 88 500 108
rect 0 48 30 88
rect 70 48 110 88
rect 150 48 190 88
rect 230 48 270 88
rect 310 48 350 88
rect 390 48 430 88
rect 470 48 500 88
rect 0 28 500 48
rect 30 -32 60 28
rect 30 -80 70 -32
rect 30 -120 40 -80
rect 30 -144 70 -120
rect 120 -80 160 -32
rect 120 -120 125 -80
rect 155 -120 160 -80
rect 120 -144 160 -120
rect 200 -80 240 -32
rect 200 -120 205 -80
rect 235 -120 240 -80
rect 200 -144 240 -120
rect 300 -80 340 -32
rect 300 -120 305 -80
rect 335 -120 340 -80
rect 300 -144 340 -120
rect 400 -80 440 -32
rect 400 -120 404 -80
rect 434 -120 440 -80
rect 400 -144 440 -120
rect 70 -190 110 -180
rect 260 -190 300 -180
rect 70 -193 300 -190
rect 70 -220 79 -193
rect 102 -194 300 -193
rect 102 -216 270 -194
rect 290 -216 300 -194
rect 102 -220 300 -216
rect 70 -230 110 -220
rect 260 -230 300 -220
rect 410 -255 440 -144
rect -10 -285 440 -255
rect 70 -324 110 -313
rect 70 -330 79 -324
rect -10 -349 79 -330
rect 102 -349 110 -324
rect -10 -360 110 -349
rect 260 -321 300 -310
rect 260 -347 268 -321
rect 294 -347 300 -321
rect 260 -360 300 -347
rect 350 -324 390 -310
rect 350 -346 360 -324
rect 380 -346 390 -324
rect 350 -360 390 -346
rect 410 -398 440 -285
rect 30 -408 70 -398
rect 30 -432 38 -408
rect 62 -432 70 -408
rect 30 -440 70 -432
rect 120 -406 160 -398
rect 120 -432 128 -406
rect 154 -432 160 -406
rect 120 -440 160 -432
rect 200 -406 240 -398
rect 200 -432 208 -406
rect 234 -432 240 -406
rect 40 -490 70 -440
rect 200 -441 240 -432
rect 300 -406 340 -398
rect 300 -432 308 -406
rect 334 -432 340 -406
rect 300 -440 340 -432
rect 400 -406 440 -398
rect 400 -432 408 -406
rect 434 -432 440 -406
rect 400 -440 440 -432
rect 0 -510 500 -490
rect 0 -550 30 -510
rect 70 -550 110 -510
rect 150 -550 190 -510
rect 230 -550 270 -510
rect 310 -550 350 -510
rect 390 -550 430 -510
rect 470 -550 500 -510
rect 0 -570 500 -550
<< viali >>
rect 125 -120 155 -80
rect 205 -120 235 -80
rect 305 -120 335 -80
rect 270 -216 290 -194
rect 268 -347 294 -321
rect 360 -346 380 -324
rect 128 -432 154 -406
rect 208 -432 234 -406
rect 308 -432 334 -406
<< metal1 >>
rect 120 -80 160 -32
rect 120 -120 125 -80
rect 155 -120 160 -80
rect 120 -144 160 -120
rect 200 -80 240 -32
rect 200 -120 205 -80
rect 235 -120 240 -80
rect 200 -144 240 -120
rect 300 -80 340 -32
rect 300 -120 305 -80
rect 335 -114 340 -80
rect 335 -120 481 -114
rect 300 -144 481 -120
rect 200 -190 230 -144
rect -10 -220 230 -190
rect 200 -398 230 -220
rect 260 -190 300 -180
rect 260 -194 380 -190
rect 260 -216 270 -194
rect 290 -216 380 -194
rect 260 -220 380 -216
rect 260 -230 300 -220
rect 350 -310 380 -220
rect 450 -255 480 -144
rect 450 -285 510 -255
rect 260 -321 300 -310
rect 260 -347 268 -321
rect 294 -347 300 -321
rect 260 -360 300 -347
rect 350 -324 390 -310
rect 350 -346 360 -324
rect 380 -346 390 -324
rect 350 -360 390 -346
rect 450 -398 480 -285
rect 120 -406 160 -398
rect 120 -432 128 -406
rect 154 -432 160 -406
rect 120 -440 160 -432
rect 200 -406 240 -398
rect 200 -432 208 -406
rect 234 -432 240 -406
rect 200 -441 240 -432
rect 300 -406 480 -398
rect 300 -432 308 -406
rect 334 -428 480 -406
rect 334 -432 340 -428
rect 300 -440 340 -432
<< via1 >>
rect 125 -120 155 -80
rect 268 -347 294 -321
rect 128 -432 154 -406
<< metal2 >>
rect 120 -80 160 -32
rect 120 -120 125 -80
rect 155 -120 160 -80
rect 120 -144 160 -120
rect 130 -320 160 -144
rect 260 -320 300 -310
rect 130 -321 300 -320
rect 130 -347 268 -321
rect 294 -347 300 -321
rect 130 -350 300 -347
rect 130 -398 160 -350
rect 260 -360 300 -350
rect 120 -406 160 -398
rect 120 -432 128 -406
rect 154 -432 160 -406
rect 120 -440 160 -432
<< labels >>
rlabel locali 240 -540 258 -530 1 gnd!
rlabel metal1 0 -210 18 -200 1 i1
rlabel locali 0 -277 18 -267 1 i2
rlabel locali 1 -350 19 -340 1 se
rlabel metal1 489 -274 507 -264 1 out
rlabel locali 241 58 259 68 1 vdd
<< end >>
