magic
tech sky130A
timestamp 1605175454
<< nwell >>
rect -75 -85 1190 379
<< nmos >>
rect 21 -670 61 -610
rect 161 -670 201 -610
rect 260 -670 300 -610
rect 374 -670 414 -610
rect 489 -670 529 -610
rect 639 -670 679 -610
rect 737 -670 777 -610
rect 894 -670 934 -610
rect 1037 -670 1077 -610
<< pmos >>
rect 21 52 61 212
rect 161 52 201 212
rect 260 52 300 212
rect 374 52 414 212
rect 489 52 529 212
rect 639 52 679 212
rect 737 52 777 212
rect 894 52 934 212
rect 1037 52 1077 212
<< ndiff >>
rect -19 -637 21 -610
rect -19 -662 -14 -637
rect 6 -662 21 -637
rect -19 -670 21 -662
rect 61 -637 96 -610
rect 61 -662 72 -637
rect 92 -662 96 -637
rect 61 -670 96 -662
rect 123 -637 161 -610
rect 123 -662 128 -637
rect 148 -662 161 -637
rect 123 -670 161 -662
rect 201 -637 260 -610
rect 201 -662 215 -637
rect 236 -662 260 -637
rect 201 -670 260 -662
rect 300 -637 374 -610
rect 300 -662 328 -637
rect 349 -662 374 -637
rect 300 -670 374 -662
rect 414 -637 489 -610
rect 414 -662 439 -637
rect 460 -662 489 -637
rect 414 -670 489 -662
rect 529 -637 572 -610
rect 529 -662 549 -637
rect 568 -662 572 -637
rect 529 -670 572 -662
rect 599 -637 639 -610
rect 599 -662 604 -637
rect 624 -662 639 -637
rect 599 -670 639 -662
rect 679 -637 737 -610
rect 679 -662 690 -637
rect 711 -662 737 -637
rect 679 -670 737 -662
rect 777 -637 826 -610
rect 777 -662 803 -637
rect 822 -662 826 -637
rect 777 -670 826 -662
rect 854 -637 894 -610
rect 854 -662 859 -637
rect 879 -662 894 -637
rect 854 -670 894 -662
rect 934 -637 969 -610
rect 934 -662 945 -637
rect 964 -662 969 -637
rect 934 -670 969 -662
rect 997 -637 1037 -610
rect 997 -662 1002 -637
rect 1022 -662 1037 -637
rect 997 -670 1037 -662
rect 1077 -637 1153 -610
rect 1077 -662 1088 -637
rect 1109 -662 1153 -637
rect 1077 -670 1153 -662
<< pdiff >>
rect -19 203 21 212
rect -19 164 -14 203
rect 6 164 21 203
rect -19 52 21 164
rect 61 173 96 212
rect 61 142 73 173
rect 92 142 96 173
rect 61 52 96 142
rect 123 203 161 212
rect 123 164 127 203
rect 147 164 161 203
rect 123 52 161 164
rect 201 173 260 212
rect 201 142 216 173
rect 235 142 260 173
rect 201 52 260 142
rect 300 173 374 212
rect 300 142 329 173
rect 348 142 374 173
rect 300 52 374 142
rect 414 173 489 212
rect 414 142 440 173
rect 459 142 489 173
rect 414 52 489 142
rect 529 173 572 212
rect 529 142 550 173
rect 568 142 572 173
rect 529 52 572 142
rect 599 203 639 212
rect 599 164 604 203
rect 624 164 639 203
rect 599 52 639 164
rect 679 173 737 212
rect 679 142 691 173
rect 710 142 737 173
rect 679 52 737 142
rect 777 173 826 212
rect 777 142 804 173
rect 822 142 826 173
rect 777 52 826 142
rect 854 203 894 212
rect 854 164 859 203
rect 879 164 894 203
rect 854 52 894 164
rect 934 173 969 212
rect 934 142 946 173
rect 965 142 969 173
rect 934 52 969 142
rect 997 203 1037 212
rect 997 164 1002 203
rect 1022 164 1037 203
rect 997 52 1037 164
rect 1077 173 1154 212
rect 1077 142 1089 173
rect 1108 142 1154 173
rect 1077 52 1154 142
<< ndiffc >>
rect -14 -662 6 -637
rect 72 -662 92 -637
rect 128 -662 148 -637
rect 215 -662 236 -637
rect 328 -662 349 -637
rect 439 -662 460 -637
rect 549 -662 568 -637
rect 604 -662 624 -637
rect 690 -662 711 -637
rect 803 -662 822 -637
rect 859 -662 879 -637
rect 945 -662 964 -637
rect 1002 -662 1022 -637
rect 1088 -662 1109 -637
<< pdiffc >>
rect -14 164 6 203
rect 73 142 92 173
rect 127 164 147 203
rect 216 142 235 173
rect 329 142 348 173
rect 440 142 459 173
rect 550 142 568 173
rect 604 164 624 203
rect 691 142 710 173
rect 804 142 822 173
rect 859 164 879 203
rect 946 142 965 173
rect 1002 164 1022 203
rect 1089 142 1108 173
<< psubdiff >>
rect -37 -744 6 -723
rect 27 -744 52 -723
rect 73 -744 1164 -723
<< nsubdiff >>
rect -40 338 535 359
rect 556 338 895 359
rect 916 338 1086 359
rect 1107 338 1170 359
<< psubdiffcont >>
rect 6 -744 27 -723
rect 52 -744 73 -723
<< nsubdiffcont >>
rect 535 338 556 359
rect 895 338 916 359
rect 1086 338 1107 359
<< poly >>
rect 21 212 61 237
rect 161 212 201 237
rect 260 212 300 237
rect 374 212 414 237
rect 489 212 529 237
rect 639 212 679 237
rect 737 212 777 237
rect 894 212 934 237
rect 1037 212 1077 237
rect 21 -375 61 52
rect 161 -313 201 52
rect 260 -85 300 52
rect 374 -28 414 52
rect 489 -28 529 52
rect 369 -38 529 -28
rect 369 -68 377 -38
rect 411 -68 529 -38
rect 369 -78 419 -68
rect 255 -95 305 -85
rect 255 -125 263 -95
rect 297 -125 305 -95
rect 255 -135 305 -125
rect 639 -149 679 52
rect 737 -85 777 52
rect 732 -95 782 -85
rect 732 -125 740 -95
rect 774 -125 782 -95
rect 732 -135 782 -125
rect 608 -159 679 -149
rect 608 -184 618 -159
rect 643 -184 679 -159
rect 608 -194 679 -184
rect 150 -323 201 -313
rect 150 -348 160 -323
rect 185 -348 201 -323
rect 150 -358 201 -348
rect -1 -385 61 -375
rect -1 -415 7 -385
rect 41 -415 61 -385
rect -1 -425 61 -415
rect 21 -610 61 -425
rect 161 -610 201 -358
rect 255 -385 305 -375
rect 255 -415 263 -385
rect 297 -415 305 -385
rect 255 -425 305 -415
rect 260 -610 300 -425
rect 479 -496 529 -486
rect 479 -526 487 -496
rect 521 -526 529 -496
rect 479 -536 529 -526
rect 374 -573 529 -536
rect 374 -610 414 -573
rect 489 -610 529 -573
rect 639 -610 679 -194
rect 894 -257 934 52
rect 1037 -149 1077 52
rect 1024 -159 1077 -149
rect 1024 -184 1034 -159
rect 1059 -184 1077 -159
rect 1024 -194 1077 -184
rect 881 -267 934 -257
rect 881 -292 891 -267
rect 916 -292 934 -267
rect 881 -302 934 -292
rect 732 -385 782 -375
rect 732 -415 740 -385
rect 774 -415 782 -385
rect 732 -425 782 -415
rect 737 -610 777 -425
rect 894 -610 934 -302
rect 1037 -610 1077 -194
rect 21 -690 61 -670
rect 161 -691 201 -670
rect 260 -691 300 -670
rect 374 -691 414 -670
rect 489 -691 529 -670
rect 639 -691 679 -670
rect 737 -691 777 -670
rect 894 -690 934 -670
rect 1037 -690 1077 -670
<< polycont >>
rect 377 -68 411 -38
rect 263 -125 297 -95
rect 740 -125 774 -95
rect 618 -184 643 -159
rect 160 -348 185 -323
rect 7 -415 41 -385
rect 263 -415 297 -385
rect 487 -526 521 -496
rect 1034 -184 1059 -159
rect 891 -292 916 -267
rect 740 -415 774 -385
<< locali >>
rect -56 359 1185 367
rect -56 338 -25 359
rect -4 338 535 359
rect 556 338 895 359
rect 916 338 1086 359
rect 1107 338 1134 359
rect 1155 338 1185 359
rect -56 332 1185 338
rect -19 203 6 332
rect -19 164 -14 203
rect -19 52 6 164
rect 70 173 96 212
rect 70 142 73 173
rect 92 142 96 173
rect 70 -206 96 142
rect 123 203 148 332
rect 123 164 127 203
rect 147 164 148 203
rect 123 52 148 164
rect 212 173 238 212
rect 212 142 216 173
rect 235 142 238 173
rect 212 -153 238 142
rect 325 173 351 212
rect 325 142 329 173
rect 348 142 351 173
rect 255 -95 305 -85
rect 255 -125 263 -95
rect 297 -125 305 -95
rect 255 -135 305 -125
rect 212 -162 249 -153
rect 212 -179 221 -162
rect 240 -179 249 -162
rect 212 -189 249 -179
rect 70 -219 120 -206
rect 70 -239 85 -219
rect 105 -239 120 -219
rect 70 -256 120 -239
rect -1 -379 49 -375
rect -25 -385 49 -379
rect -25 -409 7 -385
rect -1 -415 7 -409
rect 41 -415 49 -385
rect -1 -425 49 -415
rect -19 -637 7 -610
rect -19 -662 -14 -637
rect 6 -662 7 -637
rect -19 -715 7 -662
rect 70 -637 96 -256
rect 212 -263 238 -189
rect 212 -272 249 -263
rect 212 -289 222 -272
rect 241 -289 249 -272
rect 212 -299 249 -289
rect 150 -323 195 -313
rect 150 -348 160 -323
rect 185 -348 195 -323
rect 150 -358 195 -348
rect 70 -662 72 -637
rect 92 -662 96 -637
rect 70 -670 96 -662
rect 123 -637 149 -610
rect 123 -662 128 -637
rect 148 -662 149 -637
rect 123 -715 149 -662
rect 212 -637 238 -299
rect 255 -385 305 -375
rect 255 -415 263 -385
rect 297 -415 305 -385
rect 255 -425 305 -415
rect 212 -662 215 -637
rect 236 -662 238 -637
rect 212 -670 238 -662
rect 325 -637 351 142
rect 436 173 462 212
rect 436 142 440 173
rect 459 142 462 173
rect 369 -38 419 -28
rect 369 -68 377 -38
rect 411 -68 419 -38
rect 369 -78 419 -68
rect 436 -440 462 142
rect 546 173 572 212
rect 546 142 550 173
rect 568 142 572 173
rect 546 -315 572 142
rect 599 203 624 332
rect 599 164 604 203
rect 599 52 624 164
rect 688 173 714 212
rect 688 142 691 173
rect 710 142 714 173
rect 608 -159 653 -149
rect 608 -184 618 -159
rect 643 -184 653 -159
rect 608 -194 653 -184
rect 536 -325 573 -315
rect 536 -342 545 -325
rect 564 -342 573 -325
rect 536 -351 573 -342
rect 425 -450 462 -440
rect 425 -467 435 -450
rect 454 -467 462 -450
rect 425 -476 462 -467
rect 325 -662 328 -637
rect 349 -662 351 -637
rect 325 -670 351 -662
rect 436 -637 462 -476
rect 479 -496 529 -486
rect 479 -526 487 -496
rect 521 -526 529 -496
rect 479 -536 529 -526
rect 436 -662 439 -637
rect 460 -662 462 -637
rect 436 -670 462 -662
rect 546 -637 572 -351
rect 546 -662 549 -637
rect 568 -662 572 -637
rect 546 -670 572 -662
rect 599 -637 625 -610
rect 599 -662 604 -637
rect 624 -662 625 -637
rect 599 -715 625 -662
rect 688 -637 714 142
rect 800 173 826 212
rect 800 142 804 173
rect 822 142 826 173
rect 732 -95 782 -85
rect 732 -125 740 -95
rect 774 -125 782 -95
rect 732 -135 782 -125
rect 800 -315 826 142
rect 854 203 879 332
rect 854 164 859 203
rect 854 52 879 164
rect 943 173 969 212
rect 943 142 946 173
rect 965 142 969 173
rect 943 -153 969 142
rect 997 203 1022 332
rect 997 164 1002 203
rect 997 52 1022 164
rect 1086 173 1112 212
rect 1086 142 1089 173
rect 1108 142 1112 173
rect 943 -162 980 -153
rect 943 -179 953 -162
rect 972 -164 980 -162
rect 1024 -159 1069 -149
rect 1024 -164 1034 -159
rect 972 -179 1034 -164
rect 943 -184 1034 -179
rect 1059 -184 1069 -159
rect 943 -189 1069 -184
rect 881 -267 926 -257
rect 881 -292 891 -267
rect 916 -292 926 -267
rect 881 -302 926 -292
rect 792 -324 829 -315
rect 792 -341 802 -324
rect 821 -341 829 -324
rect 792 -351 829 -341
rect 732 -385 782 -375
rect 732 -415 740 -385
rect 774 -415 782 -385
rect 732 -425 782 -415
rect 688 -662 690 -637
rect 711 -662 714 -637
rect 688 -670 714 -662
rect 800 -637 826 -351
rect 800 -662 803 -637
rect 822 -662 826 -637
rect 800 -670 826 -662
rect 854 -637 880 -610
rect 854 -662 859 -637
rect 879 -662 880 -637
rect 854 -715 880 -662
rect 943 -637 969 -189
rect 1024 -194 1069 -189
rect 1086 -439 1112 142
rect 1085 -448 1122 -439
rect 1085 -465 1094 -448
rect 1113 -465 1122 -448
rect 1085 -475 1122 -465
rect 943 -662 945 -637
rect 964 -662 969 -637
rect 943 -670 969 -662
rect 997 -637 1023 -610
rect 997 -662 1002 -637
rect 1022 -662 1023 -637
rect 997 -715 1023 -662
rect 1086 -637 1112 -475
rect 1086 -662 1088 -637
rect 1109 -662 1112 -637
rect 1086 -670 1112 -662
rect -49 -723 1178 -715
rect -49 -744 -30 -723
rect -9 -744 6 -723
rect 27 -744 52 -723
rect 73 -744 1141 -723
rect 1162 -744 1178 -723
rect -49 -750 1178 -744
<< viali >>
rect -25 338 -4 359
rect 1134 338 1155 359
rect 263 -125 297 -95
rect 221 -179 240 -162
rect 85 -239 105 -219
rect 7 -415 41 -385
rect 222 -289 241 -272
rect 160 -348 185 -323
rect 263 -415 297 -385
rect 377 -68 411 -38
rect 618 -184 643 -159
rect 545 -342 564 -325
rect 435 -467 454 -450
rect 487 -526 521 -496
rect 740 -125 774 -95
rect 953 -179 972 -162
rect 1034 -184 1059 -159
rect 891 -292 916 -267
rect 802 -341 821 -324
rect 740 -415 774 -385
rect 1094 -465 1113 -448
rect -30 -744 -9 -723
rect 1141 -744 1162 -723
<< metal1 >>
rect -68 359 1190 371
rect -68 338 -25 359
rect -4 338 1134 359
rect 1155 338 1190 359
rect -68 327 1190 338
rect 369 -34 419 -28
rect 369 -72 374 -34
rect 414 -72 419 -34
rect 369 -78 419 -72
rect 255 -91 305 -85
rect 255 -129 260 -91
rect 300 -129 305 -91
rect 255 -135 305 -129
rect 732 -91 782 -85
rect 732 -129 737 -91
rect 777 -129 782 -91
rect 732 -135 782 -129
rect 212 -158 249 -153
rect 212 -184 218 -158
rect 244 -184 249 -158
rect 212 -189 249 -184
rect 608 -157 653 -149
rect 608 -186 616 -157
rect 645 -186 653 -157
rect 608 -194 653 -186
rect 943 -158 980 -153
rect 943 -184 949 -158
rect 975 -184 980 -158
rect 943 -189 980 -184
rect 1024 -157 1069 -149
rect 1024 -186 1032 -157
rect 1061 -186 1069 -157
rect 1024 -194 1069 -186
rect 70 -214 120 -206
rect 70 -246 80 -214
rect 112 -246 120 -214
rect 70 -256 120 -246
rect 212 -268 249 -263
rect 212 -294 218 -268
rect 244 -294 249 -268
rect 212 -299 249 -294
rect 881 -265 926 -257
rect 881 -294 889 -265
rect 918 -294 926 -265
rect 881 -302 926 -294
rect 150 -321 195 -313
rect 150 -350 158 -321
rect 187 -350 195 -321
rect 150 -358 195 -350
rect 536 -320 573 -315
rect 536 -346 542 -320
rect 568 -346 573 -320
rect 536 -351 573 -346
rect 792 -320 829 -315
rect 792 -346 798 -320
rect 824 -346 829 -320
rect 792 -351 829 -346
rect -1 -381 49 -375
rect -1 -419 4 -381
rect 44 -419 49 -381
rect -1 -425 49 -419
rect 255 -381 305 -375
rect 255 -419 260 -381
rect 300 -419 305 -381
rect 255 -425 305 -419
rect 732 -381 782 -375
rect 732 -419 737 -381
rect 777 -419 782 -381
rect 732 -425 782 -419
rect 425 -445 462 -440
rect 425 -471 431 -445
rect 457 -471 462 -445
rect 425 -476 462 -471
rect 1085 -444 1122 -439
rect 1085 -470 1091 -444
rect 1117 -470 1122 -444
rect 1085 -475 1122 -470
rect 479 -492 529 -486
rect 479 -530 484 -492
rect 524 -530 529 -492
rect 479 -536 529 -530
rect -62 -723 1193 -710
rect -62 -744 -30 -723
rect -9 -744 1141 -723
rect 1162 -744 1193 -723
rect -62 -754 1193 -744
<< via1 >>
rect 374 -38 414 -34
rect 374 -68 377 -38
rect 377 -68 411 -38
rect 411 -68 414 -38
rect 374 -72 414 -68
rect 260 -95 300 -91
rect 260 -125 263 -95
rect 263 -125 297 -95
rect 297 -125 300 -95
rect 260 -129 300 -125
rect 737 -95 777 -91
rect 737 -125 740 -95
rect 740 -125 774 -95
rect 774 -125 777 -95
rect 737 -129 777 -125
rect 218 -162 244 -158
rect 218 -179 221 -162
rect 221 -179 240 -162
rect 240 -179 244 -162
rect 218 -184 244 -179
rect 616 -159 645 -157
rect 616 -184 618 -159
rect 618 -184 643 -159
rect 643 -184 645 -159
rect 616 -186 645 -184
rect 949 -162 975 -158
rect 949 -179 953 -162
rect 953 -179 972 -162
rect 972 -179 975 -162
rect 949 -184 975 -179
rect 1032 -159 1061 -157
rect 1032 -184 1034 -159
rect 1034 -184 1059 -159
rect 1059 -184 1061 -159
rect 1032 -186 1061 -184
rect 80 -219 112 -214
rect 80 -239 85 -219
rect 85 -239 105 -219
rect 105 -239 112 -219
rect 80 -246 112 -239
rect 218 -272 244 -268
rect 218 -289 222 -272
rect 222 -289 241 -272
rect 241 -289 244 -272
rect 218 -294 244 -289
rect 889 -267 918 -265
rect 889 -292 891 -267
rect 891 -292 916 -267
rect 916 -292 918 -267
rect 889 -294 918 -292
rect 158 -323 187 -321
rect 158 -348 160 -323
rect 160 -348 185 -323
rect 185 -348 187 -323
rect 158 -350 187 -348
rect 542 -325 568 -320
rect 542 -342 545 -325
rect 545 -342 564 -325
rect 564 -342 568 -325
rect 542 -346 568 -342
rect 798 -324 824 -320
rect 798 -341 802 -324
rect 802 -341 821 -324
rect 821 -341 824 -324
rect 798 -346 824 -341
rect 4 -385 44 -381
rect 4 -415 7 -385
rect 7 -415 41 -385
rect 41 -415 44 -385
rect 4 -419 44 -415
rect 260 -385 300 -381
rect 260 -415 263 -385
rect 263 -415 297 -385
rect 297 -415 300 -385
rect 260 -419 300 -415
rect 737 -385 777 -381
rect 737 -415 740 -385
rect 740 -415 774 -385
rect 774 -415 777 -385
rect 737 -419 777 -415
rect 431 -450 457 -445
rect 431 -467 435 -450
rect 435 -467 454 -450
rect 454 -467 457 -450
rect 431 -471 457 -467
rect 1091 -448 1117 -444
rect 1091 -465 1094 -448
rect 1094 -465 1113 -448
rect 1113 -465 1117 -448
rect 1091 -470 1117 -465
rect 484 -496 524 -492
rect 484 -526 487 -496
rect 487 -526 521 -496
rect 521 -526 524 -496
rect 484 -530 524 -526
<< metal2 >>
rect 369 -34 419 -28
rect 369 -72 374 -34
rect 414 -72 419 -34
rect 369 -78 419 -72
rect 255 -91 305 -85
rect 255 -129 260 -91
rect 300 -129 305 -91
rect 255 -135 305 -129
rect 732 -91 782 -85
rect 732 -129 737 -91
rect 777 -129 782 -91
rect 732 -135 782 -129
rect 212 -158 249 -153
rect 212 -184 218 -158
rect 244 -164 249 -158
rect 608 -157 653 -149
rect 608 -164 616 -157
rect 244 -184 616 -164
rect 212 -186 616 -184
rect 645 -186 653 -157
rect 212 -189 653 -186
rect 943 -158 980 -153
rect 943 -184 949 -158
rect 975 -184 980 -158
rect 943 -189 980 -184
rect 1024 -157 1069 -149
rect 1024 -186 1032 -157
rect 1061 -164 1069 -157
rect 1061 -186 1161 -164
rect 1024 -189 1161 -186
rect 608 -194 653 -189
rect 1024 -194 1069 -189
rect 70 -214 120 -206
rect 70 -246 80 -214
rect 112 -246 120 -214
rect 70 -256 120 -246
rect 212 -268 249 -263
rect 212 -294 218 -268
rect 244 -274 249 -268
rect 881 -265 926 -257
rect 881 -274 889 -265
rect 244 -294 889 -274
rect 918 -294 926 -265
rect 212 -299 926 -294
rect 881 -302 926 -299
rect 150 -315 195 -313
rect 150 -320 829 -315
rect 150 -321 542 -320
rect 150 -350 158 -321
rect 187 -340 542 -321
rect 187 -350 195 -340
rect 150 -358 195 -350
rect 536 -346 542 -340
rect 568 -340 798 -320
rect 568 -346 573 -340
rect 536 -351 573 -346
rect 792 -346 798 -340
rect 824 -346 829 -320
rect 792 -351 829 -346
rect -1 -381 49 -375
rect -1 -419 4 -381
rect 44 -419 49 -381
rect -1 -425 49 -419
rect 255 -381 305 -375
rect 255 -419 260 -381
rect 300 -419 305 -381
rect 255 -425 305 -419
rect 732 -381 782 -375
rect 732 -419 737 -381
rect 777 -419 782 -381
rect 732 -425 782 -419
rect 1085 -440 1122 -439
rect 425 -444 1122 -440
rect 425 -445 1091 -444
rect 425 -471 431 -445
rect 457 -465 1091 -445
rect 457 -471 462 -465
rect 425 -476 462 -471
rect 1085 -470 1091 -465
rect 1117 -470 1122 -444
rect 1085 -475 1122 -470
rect 479 -492 529 -486
rect 479 -530 484 -492
rect 524 -530 529 -492
rect 479 -536 529 -530
<< via2 >>
rect 374 -72 414 -34
rect 260 -129 300 -91
rect 737 -129 777 -91
rect 80 -246 112 -214
rect 4 -419 44 -381
rect 260 -419 300 -381
rect 737 -419 777 -381
rect 484 -530 524 -492
<< metal3 >>
rect 369 -34 419 -28
rect 369 -72 374 -34
rect 414 -72 419 -34
rect 369 -78 419 -72
rect 255 -91 305 -85
rect 255 -129 260 -91
rect 300 -129 305 -91
rect 255 -135 305 -129
rect 70 -214 120 -206
rect 70 -246 80 -214
rect 112 -246 120 -214
rect 70 -256 120 -246
rect 373 -375 403 -78
rect 732 -91 782 -85
rect 732 -129 737 -91
rect 777 -129 782 -91
rect 732 -135 782 -129
rect -1 -381 782 -375
rect -1 -419 4 -381
rect 44 -405 260 -381
rect 44 -419 49 -405
rect -1 -425 49 -419
rect 255 -419 260 -405
rect 300 -405 737 -381
rect 300 -419 305 -405
rect 255 -425 305 -419
rect 732 -419 737 -405
rect 777 -419 782 -381
rect 732 -425 782 -419
rect 479 -492 529 -486
rect 479 -530 484 -492
rect 524 -530 529 -492
rect 479 -536 529 -530
<< via3 >>
rect 260 -129 300 -91
rect 80 -246 112 -214
rect 737 -129 777 -91
rect 484 -530 524 -492
<< metal4 >>
rect 255 -91 305 -85
rect 255 -129 260 -91
rect 300 -129 305 -91
rect 255 -135 305 -129
rect 732 -91 782 -85
rect 732 -129 737 -91
rect 777 -129 782 -91
rect 732 -135 782 -129
rect 257 -206 287 -135
rect 734 -206 764 -135
rect 70 -214 764 -206
rect 70 -246 80 -214
rect 112 -236 764 -214
rect 112 -246 120 -236
rect 70 -256 120 -246
rect 483 -486 513 -236
rect 479 -492 529 -486
rect 479 -530 484 -492
rect 524 -530 529 -492
rect 479 -536 529 -530
<< labels >>
flabel locali s -25 -409 -1 -379 0 FreeSans 120 0 0 0 clk
port 7 nsew
flabel metal2 s 1128 -188 1156 -165 0 FreeSans 120 0 0 0 q
port 8 nsew
flabel metal1 s 8 -735 65 -719 0 FreeSans 120 0 0 0 VGND
port 6 nsew
flabel metal1 s 30 338 95 359 0 FreeSans 120 0 0 0 VPWR
port 11 nsew
<< end >>
