
***nand1 circuit***

.include "/home/ashok/Desktop/vsd/spice_exp/sky130_fd_pr/models/corners/tt.spice"


.option scale=0.01u

Xnand in1 VDD 0 in2 out nand

.subckt nand A VPWR VGND B Y
X0 a_40_n204# A Y VGND sky130_fd_pr__nfet_01v8 w=42 l=40
X1 VPWR B Y VPWR sky130_fd_pr__pfet_01v8 w=200 l=40
X2 Y A VPWR VPWR sky130_fd_pr__pfet_01v8 w=200 l=40
X3 VGND B a_40_n204# VGND sky130_fd_pr__nfet_01v8 w=42 l=40
.ends

***set gnd and power***
 
Vdd VDD 0 1.8
Vin1 in1 0 0 pulse(0 1.8 0 10p 10p 1n 2n) 
Vin2 in2 0 0 pulse(0 1.8 0 10p 10p 0.5n 1n) 
***Vin3 in3 0 0 pulse(0 1.8 0 10p 10p 2n 4n)***
 
.op
.tran 10p 6n
.end
