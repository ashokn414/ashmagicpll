* SPICE3 file created from inv.ext - technology: sky130A

.option scale=10000u

.subckt inv A Y VPWR VGND
X0 Y A VGND VGND sky130_fd_pr__nfet_01v8 w=42 l=40
X1 Y A VPWR VPWR sky130_fd_pr__pfet_01v8 w=42 l=40
.ends
