magic
tech sky130A
timestamp 1604920739
<< nwell >>
rect -87 -62 209 139
<< nmos >>
rect 0 -204 40 -162
rect 84 -204 124 -162
<< pmos >>
rect 0 -42 40 42
rect 84 -42 124 42
<< ndiff >>
rect -40 -171 0 -162
rect -40 -196 -35 -171
rect -15 -196 0 -171
rect -40 -204 0 -196
rect 40 -204 84 -162
rect 124 -171 168 -162
rect 124 -196 143 -171
rect 163 -196 168 -171
rect 124 -204 168 -196
<< pdiff >>
rect -40 33 0 42
rect -40 -6 -35 33
rect -15 -6 0 33
rect -40 -42 0 -6
rect 40 3 84 42
rect 40 -28 52 3
rect 72 -28 84 3
rect 40 -42 84 -28
rect 124 33 168 42
rect 124 -6 143 33
rect 163 -6 168 33
rect 124 -42 168 -6
<< ndiffc >>
rect -35 -196 -15 -171
rect 143 -196 163 -171
<< pdiffc >>
rect -35 -6 -15 33
rect 52 -28 72 3
rect 143 -6 163 33
<< psubdiff >>
rect -58 -278 -15 -257
rect 6 -278 31 -257
rect 52 -278 174 -257
<< nsubdiff >>
rect -59 99 -23 120
rect -2 99 22 120
rect 43 99 174 120
<< psubdiffcont >>
rect -15 -278 6 -257
rect 31 -278 52 -257
<< nsubdiffcont >>
rect -23 99 -2 120
rect 22 99 43 120
<< poly >>
rect 0 42 40 67
rect 84 42 124 67
rect 0 -78 40 -42
rect -35 -84 40 -78
rect -35 -102 -25 -84
rect -8 -102 40 -84
rect -35 -111 40 -102
rect 0 -162 40 -111
rect 84 -78 124 -42
rect 84 -84 159 -78
rect 84 -102 132 -84
rect 149 -102 159 -84
rect 84 -111 159 -102
rect 84 -162 124 -111
rect 0 -224 40 -204
rect 84 -224 124 -204
<< polycont >>
rect -25 -102 -8 -84
rect 132 -102 149 -84
<< locali >>
rect -70 120 190 125
rect -70 99 -54 120
rect -33 99 -23 120
rect -2 99 22 120
rect 43 99 145 120
rect 166 99 190 120
rect -70 95 190 99
rect -40 33 -15 95
rect -40 -6 -35 33
rect 143 33 168 95
rect -40 -42 -15 -6
rect 49 3 75 13
rect 49 -28 52 3
rect 72 -28 75 3
rect -35 -84 0 -78
rect -35 -102 -25 -84
rect -8 -102 0 -84
rect -35 -111 0 -102
rect 49 -128 75 -28
rect 163 -6 168 33
rect 143 -42 168 -6
rect 124 -84 159 -78
rect 124 -102 132 -84
rect 149 -102 159 -84
rect 124 -111 159 -102
rect -40 -154 75 -128
rect -40 -171 -14 -154
rect -40 -196 -35 -171
rect -15 -196 -14 -171
rect -40 -204 -14 -196
rect 143 -171 168 -162
rect 163 -196 168 -171
rect 143 -249 168 -196
rect -70 -257 188 -249
rect -70 -278 -51 -257
rect -30 -278 -15 -257
rect 6 -278 31 -257
rect 52 -278 151 -257
rect 172 -278 188 -257
rect -70 -284 188 -278
<< viali >>
rect -54 99 -33 120
rect 145 99 166 120
rect -51 -278 -30 -257
rect 151 -278 172 -257
<< metal1 >>
rect -83 120 203 131
rect -83 99 -54 120
rect -33 99 145 120
rect 166 99 203 120
rect -83 88 203 99
rect -83 -257 203 -244
rect -83 -278 -51 -257
rect -30 -278 151 -257
rect 172 -278 203 -257
rect -83 -288 203 -278
<< labels >>
flabel metal1 s -10 98 56 114 0 FreeSans 120 0 0 0 VPWR
port 5 nsew
flabel locali s -25 -102 -8 -84 0 FreeSans 120 0 0 0 A
port 1 nsew
flabel metal1 s -13 -269 44 -253 0 FreeSans 120 0 0 0 VGND
port 6 nsew
flabel locali s 132 -102 149 -84 0 FreeSans 120 0 0 0 B
port 8 nsew
flabel locali s -38 -153 -18 -130 0 FreeSans 120 0 0 0 Y
port 9 nsew
<< end >>
