magic
tech sky130A
timestamp 1605695603
<< nwell >>
rect -130 -290 1245 90
rect -130 -410 1246 -290
rect -130 -1871 1263 -1491
<< nmos >>
rect 40 498 55 540
rect 200 456 215 540
rect 280 456 295 540
rect 440 498 455 540
rect 600 498 615 540
rect 760 414 775 540
rect 840 414 855 540
rect 925 414 940 540
rect 1120 498 1135 540
rect 340 -916 355 -832
rect 425 -916 440 -832
rect 600 -916 615 -832
rect 685 -916 700 -832
rect 860 -916 875 -748
rect 940 -916 955 -748
rect 1020 -916 1035 -748
rect 1100 -916 1115 -748
rect 340 -1180 355 -1096
rect 425 -1180 440 -1096
rect 600 -1180 615 -1096
rect 685 -1180 700 -1096
rect 37 -2311 52 -2269
rect 197 -2311 212 -2227
rect 277 -2311 292 -2227
rect 437 -2311 452 -2269
rect 597 -2311 612 -2269
rect 790 -2311 805 -2185
rect 870 -2311 885 -2185
rect 955 -2311 970 -2185
rect 1150 -2311 1165 -2269
<< pmos >>
rect 40 -20 55 64
rect 200 -20 215 64
rect 280 -20 295 64
rect 440 -20 455 64
rect 600 -20 615 64
rect 760 -20 775 64
rect 840 -20 855 64
rect 925 -20 940 64
rect 1120 -20 1135 64
rect 340 -384 355 -300
rect 425 -384 440 -300
rect 600 -384 615 -300
rect 685 -384 700 -300
rect 860 -384 875 -300
rect 940 -384 955 -300
rect 1020 -384 1035 -300
rect 1100 -384 1115 -300
rect 340 -1601 355 -1517
rect 425 -1601 440 -1517
rect 600 -1601 615 -1517
rect 685 -1601 700 -1517
rect 37 -1845 52 -1761
rect 197 -1845 212 -1761
rect 277 -1845 292 -1761
rect 437 -1845 452 -1761
rect 597 -1845 612 -1761
rect 790 -1845 805 -1761
rect 870 -1845 885 -1761
rect 955 -1845 970 -1761
rect 1150 -1845 1165 -1761
<< ndiff >>
rect -10 532 40 540
rect -10 508 -2 532
rect 22 508 40 532
rect -10 498 40 508
rect 55 532 110 540
rect 55 508 78 532
rect 102 508 110 532
rect 55 498 110 508
rect 150 533 200 540
rect 150 465 158 533
rect 182 465 200 533
rect 150 456 200 465
rect 215 456 280 540
rect 295 532 345 540
rect 295 464 313 532
rect 337 464 345 532
rect 390 532 440 540
rect 390 508 398 532
rect 422 508 440 532
rect 390 498 440 508
rect 455 532 510 540
rect 455 508 478 532
rect 502 508 510 532
rect 455 498 510 508
rect 550 532 600 540
rect 550 508 558 532
rect 582 508 600 532
rect 550 498 600 508
rect 615 532 670 540
rect 615 508 638 532
rect 662 508 670 532
rect 615 498 670 508
rect 710 512 760 540
rect 295 456 345 464
rect 710 444 718 512
rect 742 444 760 512
rect 710 414 760 444
rect 775 414 840 540
rect 855 414 925 540
rect 940 505 990 540
rect 940 437 958 505
rect 982 437 990 505
rect 1070 532 1120 540
rect 1070 508 1078 532
rect 1102 508 1120 532
rect 1070 498 1120 508
rect 1135 532 1190 540
rect 1135 508 1158 532
rect 1182 508 1190 532
rect 1135 498 1190 508
rect 940 414 990 437
rect 810 -780 860 -748
rect 290 -840 340 -832
rect 290 -908 298 -840
rect 322 -908 340 -840
rect 290 -916 340 -908
rect 355 -916 425 -832
rect 440 -840 490 -832
rect 440 -908 458 -840
rect 482 -908 490 -840
rect 440 -916 490 -908
rect 550 -840 600 -832
rect 550 -908 558 -840
rect 582 -908 600 -840
rect 550 -916 600 -908
rect 615 -916 685 -832
rect 700 -840 750 -832
rect 700 -908 718 -840
rect 742 -908 750 -840
rect 700 -916 750 -908
rect 810 -899 818 -780
rect 841 -899 860 -780
rect 810 -916 860 -899
rect 875 -916 940 -748
rect 955 -916 1020 -748
rect 1035 -916 1100 -748
rect 1115 -776 1171 -748
rect 1115 -897 1137 -776
rect 1163 -897 1171 -776
rect 1115 -916 1171 -897
rect 1129 -917 1171 -916
rect 450 -1096 492 -1094
rect 290 -1104 340 -1096
rect 290 -1172 298 -1104
rect 322 -1172 340 -1104
rect 290 -1180 340 -1172
rect 355 -1180 425 -1096
rect 440 -1104 492 -1096
rect 440 -1172 458 -1104
rect 484 -1172 492 -1104
rect 440 -1180 492 -1172
rect 550 -1104 600 -1096
rect 550 -1172 558 -1104
rect 582 -1172 600 -1104
rect 550 -1180 600 -1172
rect 615 -1180 685 -1096
rect 700 -1104 750 -1096
rect 700 -1172 718 -1104
rect 742 -1172 750 -1104
rect 700 -1180 750 -1172
rect 147 -2235 197 -2227
rect -13 -2279 37 -2269
rect -13 -2303 -5 -2279
rect 19 -2303 37 -2279
rect -13 -2311 37 -2303
rect 52 -2279 107 -2269
rect 52 -2303 75 -2279
rect 99 -2303 107 -2279
rect 52 -2311 107 -2303
rect 147 -2303 155 -2235
rect 179 -2303 197 -2235
rect 147 -2311 197 -2303
rect 212 -2311 277 -2227
rect 292 -2235 342 -2227
rect 292 -2303 311 -2235
rect 335 -2303 342 -2235
rect 740 -2221 790 -2185
rect 292 -2311 342 -2303
rect 387 -2279 437 -2269
rect 387 -2303 395 -2279
rect 419 -2303 437 -2279
rect 387 -2311 437 -2303
rect 452 -2279 507 -2269
rect 452 -2303 475 -2279
rect 499 -2303 507 -2279
rect 452 -2311 507 -2303
rect 547 -2279 597 -2269
rect 547 -2303 555 -2279
rect 579 -2303 597 -2279
rect 547 -2311 597 -2303
rect 612 -2279 667 -2269
rect 612 -2303 635 -2279
rect 659 -2303 667 -2279
rect 612 -2311 667 -2303
rect 740 -2289 748 -2221
rect 772 -2289 790 -2221
rect 740 -2311 790 -2289
rect 805 -2311 870 -2185
rect 885 -2311 955 -2185
rect 970 -2212 1020 -2185
rect 970 -2280 988 -2212
rect 1012 -2280 1020 -2212
rect 970 -2311 1020 -2280
rect 1100 -2279 1150 -2269
rect 1100 -2303 1108 -2279
rect 1132 -2303 1150 -2279
rect 1100 -2311 1150 -2303
rect 1165 -2279 1220 -2269
rect 1165 -2303 1188 -2279
rect 1212 -2303 1220 -2279
rect 1165 -2311 1220 -2303
<< pdiff >>
rect -10 40 40 64
rect -10 0 -4 40
rect 26 0 40 40
rect -10 -20 40 0
rect 55 40 110 64
rect 55 0 73 40
rect 103 0 110 40
rect 55 -20 110 0
rect 150 40 200 64
rect 150 0 156 40
rect 186 0 200 40
rect 150 -20 200 0
rect 215 40 280 64
rect 215 0 232 40
rect 262 0 280 40
rect 215 -20 280 0
rect 295 40 345 64
rect 295 0 310 40
rect 340 0 345 40
rect 295 -20 345 0
rect 390 40 440 64
rect 390 0 396 40
rect 426 0 440 40
rect 390 -20 440 0
rect 455 40 510 64
rect 455 0 473 40
rect 503 0 510 40
rect 455 -20 510 0
rect 550 40 600 64
rect 550 0 556 40
rect 586 0 600 40
rect 550 -20 600 0
rect 615 40 670 64
rect 615 0 633 40
rect 663 0 670 40
rect 615 -20 670 0
rect 710 40 760 64
rect 710 0 716 40
rect 746 0 760 40
rect 710 -20 760 0
rect 775 40 840 64
rect 775 0 794 40
rect 824 0 840 40
rect 775 -20 840 0
rect 855 40 925 64
rect 855 0 876 40
rect 906 0 925 40
rect 855 -20 925 0
rect 940 40 990 64
rect 940 0 955 40
rect 985 0 990 40
rect 940 -20 990 0
rect 1070 40 1120 64
rect 1070 0 1076 40
rect 1106 0 1120 40
rect 1070 -20 1120 0
rect 1135 40 1190 64
rect 1135 0 1153 40
rect 1183 0 1190 40
rect 1135 -20 1190 0
rect 290 -320 340 -300
rect 290 -360 296 -320
rect 326 -360 340 -320
rect 290 -384 340 -360
rect 355 -320 425 -300
rect 355 -360 375 -320
rect 405 -360 425 -320
rect 355 -384 425 -360
rect 440 -320 490 -300
rect 440 -360 453 -320
rect 483 -360 490 -320
rect 440 -384 490 -360
rect 550 -320 600 -300
rect 550 -360 556 -320
rect 586 -360 600 -320
rect 550 -384 600 -360
rect 615 -320 685 -300
rect 615 -360 635 -320
rect 665 -360 685 -320
rect 615 -384 685 -360
rect 700 -320 750 -300
rect 700 -360 713 -320
rect 743 -360 750 -320
rect 700 -384 750 -360
rect 810 -319 860 -300
rect 810 -359 816 -319
rect 846 -359 860 -319
rect 810 -384 860 -359
rect 875 -320 940 -300
rect 875 -360 895 -320
rect 925 -360 940 -320
rect 875 -384 940 -360
rect 955 -319 1020 -300
rect 955 -359 976 -319
rect 1006 -359 1020 -319
rect 955 -384 1020 -359
rect 1035 -319 1100 -300
rect 1035 -359 1056 -319
rect 1086 -359 1100 -319
rect 1035 -384 1100 -359
rect 1115 -319 1170 -300
rect 1115 -359 1136 -319
rect 1166 -359 1170 -319
rect 1115 -384 1170 -359
rect 290 -1541 340 -1517
rect 290 -1581 296 -1541
rect 326 -1581 340 -1541
rect 290 -1601 340 -1581
rect 355 -1541 425 -1517
rect 355 -1581 375 -1541
rect 405 -1581 425 -1541
rect 355 -1601 425 -1581
rect 440 -1541 490 -1517
rect 440 -1581 453 -1541
rect 483 -1581 490 -1541
rect 440 -1601 490 -1581
rect 550 -1541 600 -1517
rect 550 -1581 556 -1541
rect 586 -1581 600 -1541
rect 550 -1601 600 -1581
rect 615 -1541 685 -1517
rect 615 -1581 635 -1541
rect 665 -1581 685 -1541
rect 615 -1601 685 -1581
rect 700 -1541 750 -1517
rect 700 -1581 713 -1541
rect 743 -1581 750 -1541
rect 700 -1601 750 -1581
rect -13 -1781 37 -1761
rect -13 -1821 -7 -1781
rect 23 -1821 37 -1781
rect -13 -1845 37 -1821
rect 52 -1781 107 -1761
rect 52 -1821 70 -1781
rect 100 -1821 107 -1781
rect 52 -1845 107 -1821
rect 147 -1781 197 -1761
rect 147 -1821 153 -1781
rect 183 -1821 197 -1781
rect 147 -1845 197 -1821
rect 212 -1781 277 -1761
rect 212 -1821 229 -1781
rect 259 -1821 277 -1781
rect 212 -1845 277 -1821
rect 292 -1781 342 -1761
rect 292 -1821 307 -1781
rect 337 -1821 342 -1781
rect 292 -1845 342 -1821
rect 387 -1781 437 -1761
rect 387 -1821 393 -1781
rect 423 -1821 437 -1781
rect 387 -1845 437 -1821
rect 452 -1781 507 -1761
rect 452 -1821 470 -1781
rect 500 -1821 507 -1781
rect 452 -1845 507 -1821
rect 547 -1781 597 -1761
rect 547 -1821 553 -1781
rect 583 -1821 597 -1781
rect 547 -1845 597 -1821
rect 612 -1781 667 -1761
rect 612 -1821 630 -1781
rect 660 -1821 667 -1781
rect 612 -1845 667 -1821
rect 740 -1781 790 -1761
rect 740 -1821 745 -1781
rect 776 -1821 790 -1781
rect 740 -1845 790 -1821
rect 805 -1781 870 -1761
rect 805 -1821 824 -1781
rect 854 -1821 870 -1781
rect 805 -1845 870 -1821
rect 885 -1781 955 -1761
rect 885 -1821 906 -1781
rect 936 -1821 955 -1781
rect 885 -1845 955 -1821
rect 970 -1781 1020 -1761
rect 970 -1821 985 -1781
rect 1015 -1821 1020 -1781
rect 970 -1845 1020 -1821
rect 1100 -1781 1150 -1761
rect 1100 -1821 1106 -1781
rect 1136 -1821 1150 -1781
rect 1100 -1845 1150 -1821
rect 1165 -1781 1220 -1761
rect 1165 -1821 1183 -1781
rect 1213 -1821 1220 -1781
rect 1165 -1845 1220 -1821
<< ndiffc >>
rect -2 508 22 532
rect 78 508 102 532
rect 158 465 182 533
rect 313 464 337 532
rect 398 508 422 532
rect 478 508 502 532
rect 558 508 582 532
rect 638 508 662 532
rect 718 444 742 512
rect 958 437 982 505
rect 1078 508 1102 532
rect 1158 508 1182 532
rect 298 -908 322 -840
rect 458 -908 482 -840
rect 558 -908 582 -840
rect 718 -908 742 -840
rect 818 -899 841 -780
rect 1137 -897 1163 -776
rect 298 -1172 322 -1104
rect 458 -1172 484 -1104
rect 558 -1172 582 -1104
rect 718 -1172 742 -1104
rect -5 -2303 19 -2279
rect 75 -2303 99 -2279
rect 155 -2303 179 -2235
rect 311 -2303 335 -2235
rect 395 -2303 419 -2279
rect 475 -2303 499 -2279
rect 555 -2303 579 -2279
rect 635 -2303 659 -2279
rect 748 -2289 772 -2221
rect 988 -2280 1012 -2212
rect 1108 -2303 1132 -2279
rect 1188 -2303 1212 -2279
<< pdiffc >>
rect -4 0 26 40
rect 73 0 103 40
rect 156 0 186 40
rect 232 0 262 40
rect 310 0 340 40
rect 396 0 426 40
rect 473 0 503 40
rect 556 0 586 40
rect 633 0 663 40
rect 716 0 746 40
rect 794 0 824 40
rect 876 0 906 40
rect 955 0 985 40
rect 1076 0 1106 40
rect 1153 0 1183 40
rect 296 -360 326 -320
rect 375 -360 405 -320
rect 453 -360 483 -320
rect 556 -360 586 -320
rect 635 -360 665 -320
rect 713 -360 743 -320
rect 816 -359 846 -319
rect 895 -360 925 -320
rect 976 -359 1006 -319
rect 1056 -359 1086 -319
rect 1136 -359 1166 -319
rect 296 -1581 326 -1541
rect 375 -1581 405 -1541
rect 453 -1581 483 -1541
rect 556 -1581 586 -1541
rect 635 -1581 665 -1541
rect 713 -1581 743 -1541
rect -7 -1821 23 -1781
rect 70 -1821 100 -1781
rect 153 -1821 183 -1781
rect 229 -1821 259 -1781
rect 307 -1821 337 -1781
rect 393 -1821 423 -1781
rect 470 -1821 500 -1781
rect 553 -1821 583 -1781
rect 630 -1821 660 -1781
rect 745 -1821 776 -1781
rect 824 -1821 854 -1781
rect 906 -1821 936 -1781
rect 985 -1821 1015 -1781
rect 1106 -1821 1136 -1781
rect 1183 -1821 1213 -1781
<< psubdiff >>
rect -60 650 1380 660
rect -60 610 -40 650
rect 0 610 40 650
rect 80 610 120 650
rect 160 610 200 650
rect 240 610 280 650
rect 320 610 360 650
rect 400 610 440 650
rect 480 610 520 650
rect 560 610 600 650
rect 640 610 680 650
rect 720 610 760 650
rect 800 610 840 650
rect 880 610 920 650
rect 960 610 1000 650
rect 1040 610 1080 650
rect 1120 610 1160 650
rect 1200 610 1240 650
rect 1280 610 1320 650
rect 1360 610 1380 650
rect -60 600 1380 610
rect 1320 590 1380 600
rect 1320 550 1330 590
rect 1370 550 1380 590
rect 1320 510 1380 550
rect 1320 370 1330 510
rect 1370 370 1380 510
rect 1320 330 1380 370
rect 1320 290 1330 330
rect 1370 290 1380 330
rect 1320 250 1380 290
rect 1320 210 1330 250
rect 1370 210 1380 250
rect 1320 170 1380 210
rect 1320 130 1330 170
rect 1370 130 1380 170
rect 1320 90 1380 130
rect 1320 50 1330 90
rect 1370 50 1380 90
rect 1320 10 1380 50
rect 1320 -30 1330 10
rect 1370 -30 1380 10
rect 1320 -70 1380 -30
rect 1320 -170 1330 -70
rect 1370 -170 1380 -70
rect 1320 -210 1380 -170
rect 1320 -250 1330 -210
rect 1370 -250 1380 -210
rect 1320 -290 1380 -250
rect 1320 -330 1330 -290
rect 1370 -330 1380 -290
rect 1320 -370 1380 -330
rect 1320 -410 1330 -370
rect 1370 -410 1380 -370
rect 1320 -450 1380 -410
rect 1320 -490 1330 -450
rect 1370 -490 1380 -450
rect 1320 -530 1380 -490
rect 1320 -570 1330 -530
rect 1370 -570 1380 -530
rect 1320 -610 1380 -570
rect 1320 -650 1330 -610
rect 1370 -650 1380 -610
rect 1320 -690 1380 -650
rect 1320 -886 1330 -690
rect 1370 -886 1380 -690
rect 1320 -926 1380 -886
rect 1320 -966 1330 -926
rect 1370 -966 1380 -926
rect 1320 -976 1380 -966
rect 290 -986 1380 -976
rect 290 -1026 310 -986
rect 350 -1026 390 -986
rect 430 -1026 830 -986
rect 870 -1026 910 -986
rect 950 -1026 990 -986
rect 1030 -1026 1070 -986
rect 1110 -1026 1270 -986
rect 1310 -1006 1380 -986
rect 1310 -1026 1330 -1006
rect 290 -1036 1330 -1026
rect 1320 -1046 1330 -1036
rect 1370 -1046 1380 -1006
rect 1320 -1086 1380 -1046
rect 1320 -1126 1330 -1086
rect 1370 -1126 1380 -1086
rect 1320 -1211 1380 -1126
rect 1320 -1251 1330 -1211
rect 1370 -1251 1380 -1211
rect 1320 -1291 1380 -1251
rect 1320 -1331 1330 -1291
rect 1370 -1331 1380 -1291
rect 1320 -1371 1380 -1331
rect 1320 -1411 1330 -1371
rect 1370 -1411 1380 -1371
rect 1320 -1451 1380 -1411
rect 1320 -1491 1330 -1451
rect 1370 -1491 1380 -1451
rect 1320 -1531 1380 -1491
rect 1320 -1571 1330 -1531
rect 1370 -1571 1380 -1531
rect 1320 -1611 1380 -1571
rect 1320 -1651 1330 -1611
rect 1370 -1651 1380 -1611
rect 1320 -1691 1380 -1651
rect 1320 -1731 1330 -1691
rect 1370 -1731 1380 -1691
rect 1320 -1771 1380 -1731
rect 1320 -1811 1330 -1771
rect 1370 -1811 1380 -1771
rect 1320 -1851 1380 -1811
rect 1320 -1891 1330 -1851
rect 1370 -1891 1380 -1851
rect 1320 -1931 1380 -1891
rect 1320 -1971 1330 -1931
rect 1370 -1971 1380 -1931
rect 1320 -2011 1380 -1971
rect 1320 -2051 1330 -2011
rect 1370 -2051 1380 -2011
rect 1320 -2091 1380 -2051
rect 1320 -2131 1330 -2091
rect 1370 -2131 1380 -2091
rect 1320 -2261 1380 -2131
rect 1320 -2301 1330 -2261
rect 1370 -2301 1380 -2261
rect 1320 -2360 1380 -2301
rect -60 -2370 1380 -2360
rect -60 -2410 -40 -2370
rect 0 -2410 40 -2370
rect 80 -2410 120 -2370
rect 160 -2410 200 -2370
rect 240 -2410 280 -2370
rect 320 -2410 360 -2370
rect 400 -2410 440 -2370
rect 480 -2410 520 -2370
rect 560 -2410 600 -2370
rect 640 -2410 680 -2370
rect 720 -2410 760 -2370
rect 800 -2410 840 -2370
rect 880 -2410 920 -2370
rect 960 -2410 1000 -2370
rect 1040 -2410 1080 -2370
rect 1120 -2410 1160 -2370
rect 1200 -2410 1240 -2370
rect 1280 -2410 1320 -2370
rect 1360 -2410 1380 -2370
rect -60 -2420 1380 -2410
<< nsubdiff >>
rect -90 -80 1220 -70
rect -90 -120 -50 -80
rect -10 -120 20 -80
rect 60 -120 90 -80
rect 130 -120 160 -80
rect 200 -120 310 -80
rect 350 -120 740 -80
rect 780 -120 800 -80
rect 840 -120 870 -80
rect 910 -120 940 -80
rect 980 -120 1100 -80
rect 1140 -120 1160 -80
rect 1200 -120 1220 -80
rect -90 -140 1220 -120
rect -90 -180 -50 -140
rect -10 -180 20 -140
rect 60 -180 90 -140
rect 130 -180 160 -140
rect 200 -180 310 -140
rect 350 -180 740 -140
rect 780 -180 800 -140
rect 840 -180 870 -140
rect 910 -180 940 -140
rect 980 -180 1100 -140
rect 1140 -180 1160 -140
rect 1200 -180 1220 -140
rect -90 -190 1220 -180
rect -90 -1661 1230 -1651
rect -90 -1701 -70 -1661
rect -30 -1701 0 -1661
rect 40 -1701 70 -1661
rect 110 -1701 140 -1661
rect 180 -1701 300 -1661
rect 340 -1701 750 -1661
rect 790 -1701 820 -1661
rect 860 -1701 890 -1661
rect 930 -1701 960 -1661
rect 1000 -1701 1100 -1661
rect 1140 -1701 1170 -1661
rect 1210 -1701 1230 -1661
rect -90 -1711 1230 -1701
<< psubdiffcont >>
rect -40 610 0 650
rect 40 610 80 650
rect 120 610 160 650
rect 200 610 240 650
rect 280 610 320 650
rect 360 610 400 650
rect 440 610 480 650
rect 520 610 560 650
rect 600 610 640 650
rect 680 610 720 650
rect 760 610 800 650
rect 840 610 880 650
rect 920 610 960 650
rect 1000 610 1040 650
rect 1080 610 1120 650
rect 1160 610 1200 650
rect 1240 610 1280 650
rect 1320 610 1360 650
rect 1330 550 1370 590
rect 1330 370 1370 510
rect 1330 290 1370 330
rect 1330 210 1370 250
rect 1330 130 1370 170
rect 1330 50 1370 90
rect 1330 -30 1370 10
rect 1330 -170 1370 -70
rect 1330 -250 1370 -210
rect 1330 -330 1370 -290
rect 1330 -410 1370 -370
rect 1330 -490 1370 -450
rect 1330 -570 1370 -530
rect 1330 -650 1370 -610
rect 1330 -886 1370 -690
rect 1330 -966 1370 -926
rect 310 -1026 350 -986
rect 390 -1026 430 -986
rect 830 -1026 870 -986
rect 910 -1026 950 -986
rect 990 -1026 1030 -986
rect 1070 -1026 1110 -986
rect 1270 -1026 1310 -986
rect 1330 -1046 1370 -1006
rect 1330 -1126 1370 -1086
rect 1330 -1251 1370 -1211
rect 1330 -1331 1370 -1291
rect 1330 -1411 1370 -1371
rect 1330 -1491 1370 -1451
rect 1330 -1571 1370 -1531
rect 1330 -1651 1370 -1611
rect 1330 -1731 1370 -1691
rect 1330 -1811 1370 -1771
rect 1330 -1891 1370 -1851
rect 1330 -1971 1370 -1931
rect 1330 -2051 1370 -2011
rect 1330 -2131 1370 -2091
rect 1330 -2301 1370 -2261
rect -40 -2410 0 -2370
rect 40 -2410 80 -2370
rect 120 -2410 160 -2370
rect 200 -2410 240 -2370
rect 280 -2410 320 -2370
rect 360 -2410 400 -2370
rect 440 -2410 480 -2370
rect 520 -2410 560 -2370
rect 600 -2410 640 -2370
rect 680 -2410 720 -2370
rect 760 -2410 800 -2370
rect 840 -2410 880 -2370
rect 920 -2410 960 -2370
rect 1000 -2410 1040 -2370
rect 1080 -2410 1120 -2370
rect 1160 -2410 1200 -2370
rect 1240 -2410 1280 -2370
rect 1320 -2410 1360 -2370
<< nsubdiffcont >>
rect -50 -120 -10 -80
rect 20 -120 60 -80
rect 90 -120 130 -80
rect 160 -120 200 -80
rect 310 -120 350 -80
rect 740 -120 780 -80
rect 800 -120 840 -80
rect 870 -120 910 -80
rect 940 -120 980 -80
rect 1100 -120 1140 -80
rect 1160 -120 1200 -80
rect -50 -180 -10 -140
rect 20 -180 60 -140
rect 90 -180 130 -140
rect 160 -180 200 -140
rect 310 -180 350 -140
rect 740 -180 780 -140
rect 800 -180 840 -140
rect 870 -180 910 -140
rect 940 -180 980 -140
rect 1100 -180 1140 -140
rect 1160 -180 1200 -140
rect -70 -1701 -30 -1661
rect 0 -1701 40 -1661
rect 70 -1701 110 -1661
rect 140 -1701 180 -1661
rect 300 -1701 340 -1661
rect 750 -1701 790 -1661
rect 820 -1701 860 -1661
rect 890 -1701 930 -1661
rect 960 -1701 1000 -1661
rect 1100 -1701 1140 -1661
rect 1170 -1701 1210 -1661
<< poly >>
rect 40 540 55 560
rect 200 540 215 560
rect 280 540 295 560
rect 440 540 455 560
rect 600 540 615 560
rect 760 540 775 560
rect 840 540 855 560
rect 925 540 940 560
rect 1120 540 1135 560
rect 40 240 55 498
rect 200 380 215 456
rect 175 370 215 380
rect 175 350 185 370
rect 205 350 215 370
rect 175 340 215 350
rect 15 230 55 240
rect 15 210 25 230
rect 45 210 55 230
rect 15 200 55 210
rect 40 64 55 200
rect 200 64 215 340
rect 280 333 295 456
rect 252 324 295 333
rect 252 297 261 324
rect 287 297 295 324
rect 252 290 295 297
rect 280 140 295 290
rect 440 191 455 498
rect 600 250 615 498
rect 570 240 615 250
rect 570 220 580 240
rect 600 220 615 240
rect 570 210 615 220
rect 410 181 455 191
rect 410 161 420 181
rect 440 161 455 181
rect 410 151 455 161
rect 280 130 320 140
rect 280 110 290 130
rect 310 110 320 130
rect 280 100 320 110
rect 280 64 295 100
rect 440 64 455 151
rect 600 64 615 210
rect 760 200 775 414
rect 840 283 855 414
rect 812 274 855 283
rect 812 247 821 274
rect 847 247 855 274
rect 812 240 855 247
rect 730 190 775 200
rect 730 170 740 190
rect 760 170 775 190
rect 730 160 775 170
rect 760 64 775 160
rect 840 64 855 240
rect 925 243 940 414
rect 1120 370 1135 498
rect 1095 360 1135 370
rect 1095 340 1105 360
rect 1125 340 1135 360
rect 1095 330 1135 340
rect 925 234 968 243
rect 925 207 934 234
rect 960 207 968 234
rect 925 200 968 207
rect 925 64 940 200
rect 1120 64 1135 330
rect 40 -40 55 -20
rect 200 -40 215 -20
rect 280 -40 295 -20
rect 440 -40 455 -20
rect 600 -40 615 -20
rect 760 -40 775 -20
rect 840 -40 855 -20
rect 925 -40 940 -20
rect 1120 -40 1135 -20
rect 340 -300 355 -280
rect 425 -300 440 -280
rect 600 -300 615 -280
rect 685 -300 700 -280
rect 860 -300 875 -280
rect 940 -300 955 -280
rect 1020 -300 1035 -280
rect 1100 -300 1115 -280
rect 340 -510 355 -384
rect 310 -524 355 -510
rect 310 -550 320 -524
rect 346 -550 355 -524
rect 310 -560 355 -550
rect 340 -832 355 -560
rect 425 -420 440 -384
rect 425 -430 465 -420
rect 425 -450 434 -430
rect 456 -450 465 -430
rect 425 -460 465 -450
rect 425 -832 440 -460
rect 600 -570 615 -384
rect 575 -580 615 -570
rect 575 -600 584 -580
rect 606 -600 615 -580
rect 575 -610 615 -600
rect 600 -832 615 -610
rect 685 -410 700 -384
rect 685 -420 725 -410
rect 685 -440 694 -420
rect 716 -440 725 -420
rect 685 -450 725 -440
rect 685 -832 700 -450
rect 860 -570 875 -384
rect 835 -580 875 -570
rect 835 -600 844 -580
rect 866 -600 875 -580
rect 835 -610 875 -600
rect 860 -748 875 -610
rect 940 -630 955 -384
rect 1020 -510 1035 -384
rect 990 -524 1035 -510
rect 990 -550 1000 -524
rect 1026 -550 1035 -524
rect 990 -560 1035 -550
rect 910 -644 955 -630
rect 910 -670 920 -644
rect 946 -670 955 -644
rect 910 -680 955 -670
rect 940 -748 955 -680
rect 1020 -748 1035 -560
rect 1100 -630 1115 -384
rect 1070 -644 1115 -630
rect 1070 -670 1080 -644
rect 1106 -670 1115 -644
rect 1070 -680 1115 -670
rect 1100 -748 1115 -680
rect 340 -936 355 -916
rect 425 -936 440 -916
rect 600 -936 615 -916
rect 685 -936 700 -916
rect 860 -936 875 -916
rect 940 -936 955 -916
rect 1020 -936 1035 -916
rect 1100 -936 1115 -916
rect 340 -1096 355 -1076
rect 425 -1096 440 -1076
rect 600 -1096 615 -1076
rect 685 -1096 700 -1076
rect 340 -1231 355 -1180
rect 310 -1241 355 -1231
rect 310 -1267 320 -1241
rect 346 -1267 355 -1241
rect 310 -1281 355 -1267
rect 340 -1341 355 -1281
rect 310 -1351 355 -1341
rect 310 -1377 320 -1351
rect 346 -1377 355 -1351
rect 310 -1391 355 -1377
rect 340 -1517 355 -1391
rect 425 -1441 440 -1180
rect 600 -1371 615 -1180
rect 575 -1381 615 -1371
rect 575 -1401 584 -1381
rect 606 -1401 615 -1381
rect 575 -1411 615 -1401
rect 425 -1451 465 -1441
rect 425 -1471 434 -1451
rect 456 -1471 465 -1451
rect 425 -1481 465 -1471
rect 425 -1517 440 -1481
rect 600 -1517 615 -1411
rect 685 -1301 700 -1180
rect 685 -1311 725 -1301
rect 685 -1331 694 -1311
rect 716 -1331 725 -1311
rect 685 -1341 725 -1331
rect 685 -1517 700 -1341
rect 340 -1621 355 -1601
rect 425 -1621 440 -1601
rect 600 -1621 615 -1601
rect 685 -1621 700 -1601
rect 37 -1761 52 -1741
rect 197 -1761 212 -1741
rect 277 -1761 292 -1741
rect 437 -1761 452 -1741
rect 597 -1761 612 -1741
rect 790 -1761 805 -1741
rect 870 -1761 885 -1741
rect 955 -1761 970 -1741
rect 1150 -1761 1165 -1741
rect 37 -1981 52 -1845
rect 12 -1991 52 -1981
rect 12 -2011 22 -1991
rect 42 -2011 52 -1991
rect 12 -2021 52 -2011
rect 37 -2269 52 -2021
rect 197 -2121 212 -1845
rect 277 -1881 292 -1845
rect 277 -1891 317 -1881
rect 277 -1911 287 -1891
rect 307 -1911 317 -1891
rect 277 -1921 317 -1911
rect 277 -2071 292 -1921
rect 437 -1932 452 -1845
rect 407 -1942 452 -1932
rect 407 -1962 417 -1942
rect 437 -1962 452 -1942
rect 407 -1972 452 -1962
rect 249 -2078 292 -2071
rect 249 -2105 258 -2078
rect 284 -2105 292 -2078
rect 249 -2114 292 -2105
rect 172 -2131 212 -2121
rect 172 -2151 182 -2131
rect 202 -2151 212 -2131
rect 172 -2161 212 -2151
rect 197 -2227 212 -2161
rect 277 -2227 292 -2114
rect 437 -2269 452 -1972
rect 597 -1991 612 -1845
rect 790 -1941 805 -1845
rect 760 -1951 805 -1941
rect 760 -1971 770 -1951
rect 790 -1971 805 -1951
rect 760 -1981 805 -1971
rect 567 -2001 612 -1991
rect 567 -2021 577 -2001
rect 597 -2021 612 -2001
rect 567 -2031 612 -2021
rect 597 -2269 612 -2031
rect 790 -2185 805 -1981
rect 870 -2021 885 -1845
rect 842 -2028 885 -2021
rect 842 -2055 851 -2028
rect 877 -2055 885 -2028
rect 842 -2064 885 -2055
rect 870 -2185 885 -2064
rect 955 -1981 970 -1845
rect 955 -1988 998 -1981
rect 955 -2015 964 -1988
rect 990 -2015 998 -1988
rect 955 -2024 998 -2015
rect 955 -2185 970 -2024
rect 1150 -2111 1165 -1845
rect 1125 -2121 1165 -2111
rect 1125 -2141 1135 -2121
rect 1155 -2141 1165 -2121
rect 1125 -2151 1165 -2141
rect 1150 -2269 1165 -2151
rect 37 -2331 52 -2311
rect 197 -2331 212 -2311
rect 277 -2331 292 -2311
rect 437 -2331 452 -2311
rect 597 -2331 612 -2311
rect 790 -2331 805 -2311
rect 870 -2331 885 -2311
rect 955 -2331 970 -2311
rect 1150 -2331 1165 -2311
<< polycont >>
rect 185 350 205 370
rect 25 210 45 230
rect 261 297 287 324
rect 580 220 600 240
rect 420 161 440 181
rect 290 110 310 130
rect 821 247 847 274
rect 740 170 760 190
rect 1105 340 1125 360
rect 934 207 960 234
rect 320 -550 346 -524
rect 434 -450 456 -430
rect 584 -600 606 -580
rect 694 -440 716 -420
rect 844 -600 866 -580
rect 1000 -550 1026 -524
rect 920 -670 946 -644
rect 1080 -670 1106 -644
rect 320 -1267 346 -1241
rect 320 -1377 346 -1351
rect 584 -1401 606 -1381
rect 434 -1471 456 -1451
rect 694 -1331 716 -1311
rect 22 -2011 42 -1991
rect 287 -1911 307 -1891
rect 417 -1962 437 -1942
rect 258 -2105 284 -2078
rect 182 -2151 202 -2131
rect 770 -1971 790 -1951
rect 577 -2021 597 -2001
rect 851 -2055 877 -2028
rect 964 -2015 990 -1988
rect 1135 -2141 1155 -2121
<< locali >>
rect -70 650 1390 670
rect -70 610 -40 650
rect 0 610 40 650
rect 80 610 120 650
rect 160 610 200 650
rect 240 610 280 650
rect 320 610 360 650
rect 400 610 440 650
rect 480 610 520 650
rect 560 610 600 650
rect 640 610 680 650
rect 720 610 760 650
rect 800 610 840 650
rect 880 610 920 650
rect 960 610 1000 650
rect 1040 610 1080 650
rect 1120 610 1160 650
rect 1200 610 1240 650
rect 1280 610 1320 650
rect 1360 610 1390 650
rect -70 590 1390 610
rect -10 540 20 590
rect 150 540 180 590
rect 390 540 420 590
rect 550 540 580 590
rect 710 540 740 590
rect 1070 540 1100 590
rect 1310 550 1330 590
rect 1370 550 1390 590
rect -10 532 30 540
rect -10 508 -2 532
rect 22 508 30 532
rect -10 498 30 508
rect 70 532 110 540
rect 70 508 78 532
rect 102 508 110 532
rect 70 498 110 508
rect 80 370 110 498
rect 150 533 190 540
rect 150 465 158 533
rect 182 465 190 533
rect 150 456 190 465
rect 305 532 345 540
rect 305 464 313 532
rect 337 464 345 532
rect 390 532 430 540
rect 390 508 398 532
rect 422 508 430 532
rect 390 498 430 508
rect 470 532 510 540
rect 470 508 478 532
rect 502 508 510 532
rect 470 498 510 508
rect 550 532 590 540
rect 550 508 558 532
rect 582 508 590 532
rect 550 498 590 508
rect 630 532 670 540
rect 630 508 638 532
rect 662 508 670 532
rect 630 498 670 508
rect 305 456 345 464
rect 175 370 215 380
rect 80 350 185 370
rect 205 350 215 370
rect 80 340 215 350
rect 15 230 55 240
rect -30 210 25 230
rect 45 210 55 230
rect -30 200 55 210
rect 80 64 110 340
rect 252 324 295 333
rect 252 297 261 324
rect 287 297 295 324
rect 252 290 295 297
rect 315 191 345 456
rect 480 240 510 498
rect 570 240 610 250
rect 480 220 580 240
rect 600 220 610 240
rect 480 210 610 220
rect 231 181 450 191
rect 231 161 420 181
rect 440 161 450 181
rect 231 64 261 161
rect 410 151 450 161
rect 280 130 320 140
rect 280 110 290 130
rect 310 110 320 130
rect 280 100 320 110
rect 480 64 510 210
rect 640 190 670 498
rect 710 512 750 540
rect 710 444 718 512
rect 742 444 750 512
rect 710 414 750 444
rect 950 505 990 540
rect 950 437 958 505
rect 982 437 990 505
rect 1070 532 1110 540
rect 1070 508 1078 532
rect 1102 508 1110 532
rect 1070 498 1110 508
rect 1150 532 1190 540
rect 1150 508 1158 532
rect 1182 508 1190 532
rect 1150 498 1190 508
rect 950 414 990 437
rect 950 370 980 414
rect 874 360 1135 370
rect 874 340 1105 360
rect 1125 340 1135 360
rect 700 333 740 340
rect 700 307 707 333
rect 733 330 740 333
rect 874 330 904 340
rect 1095 330 1135 340
rect 733 307 904 330
rect 700 300 904 307
rect 812 274 855 283
rect 812 247 821 274
rect 847 247 855 274
rect 812 240 855 247
rect 730 190 770 200
rect 640 170 740 190
rect 760 170 770 190
rect 640 160 770 170
rect 640 64 670 160
rect 790 130 830 140
rect 874 130 904 300
rect 925 234 968 243
rect 925 207 934 234
rect 960 207 968 234
rect 925 200 968 207
rect 1160 180 1190 498
rect 1310 510 1390 550
rect 1310 370 1330 510
rect 1370 370 1390 510
rect 1310 330 1390 370
rect 1310 290 1330 330
rect 1370 290 1390 330
rect 1310 250 1390 290
rect 1310 210 1330 250
rect 1370 210 1390 250
rect 1160 150 1230 180
rect 1310 170 1390 210
rect 790 110 800 130
rect 820 110 990 130
rect 790 100 990 110
rect 793 64 823 100
rect 960 64 990 100
rect 1160 64 1190 150
rect -10 40 30 64
rect -10 0 -4 40
rect 26 0 30 40
rect -10 -20 30 0
rect 70 40 110 64
rect 70 0 73 40
rect 103 0 110 40
rect 70 -20 110 0
rect 150 40 190 64
rect 150 0 156 40
rect 186 0 190 40
rect 150 -20 190 0
rect 227 40 267 64
rect 227 0 232 40
rect 262 0 267 40
rect 227 -20 267 0
rect 305 40 345 64
rect 305 0 310 40
rect 340 0 345 40
rect 305 -20 345 0
rect -10 -60 20 -20
rect 150 -60 180 -20
rect 315 -60 345 -20
rect 390 40 430 64
rect 390 0 396 40
rect 426 0 430 40
rect 390 -20 430 0
rect 470 40 510 64
rect 470 0 473 40
rect 503 0 510 40
rect 470 -20 510 0
rect 550 40 590 64
rect 550 0 556 40
rect 586 0 590 40
rect 550 -20 590 0
rect 630 40 670 64
rect 630 0 633 40
rect 663 0 670 40
rect 630 -20 670 0
rect 710 40 750 64
rect 710 0 716 40
rect 746 0 750 40
rect 710 -20 750 0
rect 788 40 828 64
rect 788 0 794 40
rect 824 0 828 40
rect 788 -20 828 0
rect 870 40 910 64
rect 870 0 876 40
rect 906 0 910 40
rect 870 -20 910 0
rect 950 40 990 64
rect 950 0 955 40
rect 985 0 990 40
rect 950 -20 990 0
rect 1070 40 1110 64
rect 1070 0 1076 40
rect 1106 0 1110 40
rect 1070 -20 1110 0
rect 1150 40 1190 64
rect 1150 0 1153 40
rect 1183 0 1190 40
rect 1150 -20 1190 0
rect 1310 130 1330 170
rect 1370 130 1390 170
rect 1310 90 1390 130
rect 1310 50 1330 90
rect 1370 50 1390 90
rect 1310 10 1390 50
rect 390 -60 420 -20
rect 550 -60 580 -20
rect 710 -60 740 -20
rect 870 -60 900 -20
rect 1070 -60 1100 -20
rect 1310 -30 1330 10
rect 1370 -30 1390 10
rect -130 -80 1245 -60
rect -130 -120 -50 -80
rect -10 -120 20 -80
rect 60 -120 90 -80
rect 130 -120 160 -80
rect 200 -120 310 -80
rect 350 -120 740 -80
rect 780 -120 800 -80
rect 840 -120 870 -80
rect 910 -120 940 -80
rect 980 -120 1100 -80
rect 1140 -120 1160 -80
rect 1200 -120 1245 -80
rect -130 -140 1245 -120
rect -130 -180 -50 -140
rect -10 -180 20 -140
rect 60 -180 90 -140
rect 130 -180 160 -140
rect 200 -180 310 -140
rect 350 -180 740 -140
rect 780 -180 800 -140
rect 840 -180 870 -140
rect 910 -180 940 -140
rect 980 -180 1100 -140
rect 1140 -180 1160 -140
rect 1200 -180 1245 -140
rect -130 -200 1245 -180
rect 1310 -70 1390 -30
rect 1310 -170 1330 -70
rect 1370 -170 1390 -70
rect -130 -1641 -50 -200
rect 290 -300 320 -200
rect 460 -300 490 -200
rect 290 -320 330 -300
rect 290 -360 296 -320
rect 326 -360 330 -320
rect 290 -384 330 -360
rect 370 -320 410 -300
rect 370 -360 375 -320
rect 405 -360 410 -320
rect 370 -384 410 -360
rect 450 -320 490 -300
rect 450 -360 453 -320
rect 483 -360 490 -320
rect 450 -384 490 -360
rect 550 -300 580 -200
rect 720 -300 750 -200
rect 550 -320 590 -300
rect 550 -360 556 -320
rect 586 -360 590 -320
rect 550 -384 590 -360
rect 630 -320 670 -300
rect 630 -360 635 -320
rect 665 -360 670 -320
rect 630 -384 670 -360
rect 710 -320 750 -300
rect 710 -360 713 -320
rect 743 -360 750 -320
rect 710 -384 750 -360
rect 810 -300 840 -200
rect 970 -300 1000 -200
rect 1130 -300 1160 -200
rect 1310 -210 1390 -170
rect 1310 -250 1330 -210
rect 1370 -250 1390 -210
rect 1310 -290 1390 -250
rect 810 -319 850 -300
rect 810 -359 816 -319
rect 846 -359 850 -319
rect 810 -384 850 -359
rect 890 -320 930 -300
rect 890 -360 895 -320
rect 925 -360 930 -320
rect 890 -384 930 -360
rect 970 -319 1010 -300
rect 970 -359 976 -319
rect 1006 -359 1010 -319
rect 970 -384 1010 -359
rect 1050 -319 1090 -300
rect 1050 -359 1056 -319
rect 1086 -359 1090 -319
rect 1050 -384 1090 -359
rect 1130 -319 1170 -300
rect 1130 -359 1136 -319
rect 1166 -359 1170 -319
rect 1130 -384 1170 -359
rect 1310 -330 1330 -290
rect 1370 -330 1390 -290
rect 1310 -370 1390 -330
rect 374 -480 404 -384
rect 634 -420 664 -384
rect 425 -430 664 -420
rect 425 -450 434 -430
rect 456 -450 664 -430
rect 685 -420 725 -410
rect 890 -420 920 -384
rect 1060 -420 1090 -384
rect 685 -440 694 -420
rect 716 -440 1090 -420
rect 685 -450 1090 -440
rect 425 -460 465 -450
rect 634 -470 664 -450
rect 374 -510 490 -480
rect 634 -500 750 -470
rect 310 -524 355 -510
rect 310 -550 320 -524
rect 346 -550 355 -524
rect 310 -560 355 -550
rect 460 -580 490 -510
rect 575 -580 615 -570
rect 460 -600 584 -580
rect 606 -600 615 -580
rect 460 -610 615 -600
rect 460 -832 490 -610
rect 720 -832 750 -500
rect 990 -524 1035 -510
rect 990 -550 1000 -524
rect 1026 -550 1035 -524
rect 990 -560 1035 -550
rect 1060 -560 1090 -450
rect 1310 -410 1330 -370
rect 1370 -410 1390 -370
rect 1310 -450 1390 -410
rect 1310 -490 1330 -450
rect 1370 -490 1390 -450
rect 1310 -530 1390 -490
rect 835 -580 875 -570
rect 835 -600 844 -580
rect 866 -600 875 -580
rect 1060 -590 1170 -560
rect 835 -610 875 -600
rect 910 -644 955 -630
rect 910 -670 920 -644
rect 946 -670 955 -644
rect 910 -680 955 -670
rect 1070 -644 1115 -630
rect 1070 -670 1080 -644
rect 1106 -670 1115 -644
rect 1070 -680 1115 -670
rect 1140 -748 1170 -590
rect 1310 -570 1330 -530
rect 1370 -570 1390 -530
rect 1310 -610 1390 -570
rect 1310 -650 1330 -610
rect 1370 -650 1390 -610
rect 1310 -690 1390 -650
rect 290 -840 330 -832
rect 290 -908 298 -840
rect 322 -908 330 -840
rect 290 -916 330 -908
rect 450 -840 490 -832
rect 450 -908 458 -840
rect 482 -908 490 -840
rect 450 -916 490 -908
rect 550 -840 590 -832
rect 550 -908 558 -840
rect 582 -908 590 -840
rect 550 -916 590 -908
rect 710 -840 750 -832
rect 710 -908 718 -840
rect 742 -908 750 -840
rect 710 -916 750 -908
rect 810 -780 850 -748
rect 810 -899 818 -780
rect 841 -899 850 -780
rect 810 -916 850 -899
rect 1129 -776 1171 -748
rect 1129 -897 1137 -776
rect 1163 -897 1171 -776
rect 290 -966 320 -916
rect 550 -966 580 -916
rect 810 -966 840 -916
rect 1129 -917 1171 -897
rect 1310 -886 1330 -690
rect 1370 -886 1390 -690
rect 1310 -926 1390 -886
rect 1310 -966 1330 -926
rect 1370 -966 1390 -926
rect 280 -986 1390 -966
rect 280 -1026 310 -986
rect 350 -1026 390 -986
rect 430 -1026 830 -986
rect 870 -1026 910 -986
rect 950 -1026 990 -986
rect 1030 -1026 1070 -986
rect 1110 -1026 1270 -986
rect 1310 -1006 1390 -986
rect 1310 -1026 1330 -1006
rect 280 -1046 1330 -1026
rect 1370 -1046 1390 -1006
rect 290 -1096 320 -1046
rect 290 -1104 330 -1096
rect 290 -1172 298 -1104
rect 322 -1172 330 -1104
rect 290 -1180 330 -1172
rect 450 -1104 492 -1094
rect 450 -1172 458 -1104
rect 484 -1172 492 -1104
rect 450 -1180 492 -1172
rect 550 -1096 580 -1046
rect 1310 -1086 1390 -1046
rect 550 -1104 590 -1096
rect 550 -1172 558 -1104
rect 582 -1172 590 -1104
rect 550 -1180 590 -1172
rect 710 -1104 750 -1096
rect 710 -1172 718 -1104
rect 742 -1172 750 -1104
rect 1128 -1112 1170 -1105
rect 1128 -1138 1136 -1112
rect 1162 -1138 1170 -1112
rect 1128 -1146 1170 -1138
rect 710 -1180 750 -1172
rect 310 -1241 355 -1231
rect 310 -1267 320 -1241
rect 346 -1267 355 -1241
rect 310 -1281 355 -1267
rect 310 -1351 355 -1341
rect 310 -1377 320 -1351
rect 346 -1377 355 -1351
rect 460 -1371 490 -1180
rect 720 -1201 750 -1180
rect 634 -1231 750 -1201
rect 310 -1391 355 -1377
rect 374 -1381 615 -1371
rect 374 -1401 584 -1381
rect 606 -1401 615 -1381
rect 374 -1517 404 -1401
rect 575 -1411 615 -1401
rect 425 -1451 465 -1441
rect 634 -1451 664 -1231
rect 1140 -1301 1170 -1146
rect 685 -1311 1170 -1301
rect 685 -1331 694 -1311
rect 716 -1331 1170 -1311
rect 1310 -1126 1330 -1086
rect 1370 -1126 1390 -1086
rect 1310 -1211 1390 -1126
rect 1310 -1251 1330 -1211
rect 1370 -1251 1390 -1211
rect 1310 -1291 1390 -1251
rect 1310 -1331 1330 -1291
rect 1370 -1331 1390 -1291
rect 685 -1341 725 -1331
rect 1053 -1420 1083 -1331
rect 1310 -1371 1390 -1331
rect 1310 -1411 1330 -1371
rect 1370 -1411 1390 -1371
rect 425 -1471 434 -1451
rect 456 -1471 664 -1451
rect 1043 -1427 1085 -1420
rect 1043 -1453 1051 -1427
rect 1077 -1453 1085 -1427
rect 1043 -1461 1085 -1453
rect 1310 -1451 1390 -1411
rect 425 -1481 664 -1471
rect 634 -1517 664 -1481
rect 1310 -1491 1330 -1451
rect 1370 -1491 1390 -1451
rect 290 -1541 330 -1517
rect 290 -1581 296 -1541
rect 326 -1581 330 -1541
rect 290 -1601 330 -1581
rect 370 -1541 410 -1517
rect 370 -1581 375 -1541
rect 405 -1581 410 -1541
rect 370 -1601 410 -1581
rect 450 -1541 490 -1517
rect 450 -1581 453 -1541
rect 483 -1581 490 -1541
rect 450 -1601 490 -1581
rect 290 -1641 320 -1601
rect 460 -1641 490 -1601
rect 550 -1541 590 -1517
rect 550 -1581 556 -1541
rect 586 -1581 590 -1541
rect 550 -1601 590 -1581
rect 630 -1541 670 -1517
rect 630 -1581 635 -1541
rect 665 -1581 670 -1541
rect 630 -1601 670 -1581
rect 710 -1541 750 -1517
rect 710 -1581 713 -1541
rect 743 -1581 750 -1541
rect 710 -1601 750 -1581
rect 550 -1641 580 -1601
rect 720 -1641 750 -1601
rect 1310 -1531 1390 -1491
rect 1310 -1571 1330 -1531
rect 1370 -1571 1390 -1531
rect 1310 -1611 1390 -1571
rect -130 -1661 1250 -1641
rect -130 -1701 -70 -1661
rect -30 -1701 0 -1661
rect 40 -1701 70 -1661
rect 110 -1701 140 -1661
rect 180 -1701 300 -1661
rect 340 -1701 750 -1661
rect 790 -1701 820 -1661
rect 860 -1701 890 -1661
rect 930 -1701 960 -1661
rect 1000 -1701 1100 -1661
rect 1140 -1701 1170 -1661
rect 1210 -1701 1250 -1661
rect -130 -1721 1250 -1701
rect 1310 -1651 1330 -1611
rect 1370 -1651 1390 -1611
rect 1310 -1691 1390 -1651
rect -13 -1761 17 -1721
rect 147 -1761 177 -1721
rect 312 -1761 342 -1721
rect -13 -1781 27 -1761
rect -13 -1821 -7 -1781
rect 23 -1821 27 -1781
rect -13 -1845 27 -1821
rect 67 -1781 107 -1761
rect 67 -1821 70 -1781
rect 100 -1821 107 -1781
rect 67 -1845 107 -1821
rect 147 -1781 187 -1761
rect 147 -1821 153 -1781
rect 183 -1821 187 -1781
rect 147 -1845 187 -1821
rect 224 -1781 264 -1761
rect 224 -1821 229 -1781
rect 259 -1821 264 -1781
rect 224 -1845 264 -1821
rect 302 -1781 342 -1761
rect 302 -1821 307 -1781
rect 337 -1821 342 -1781
rect 302 -1845 342 -1821
rect 387 -1761 417 -1721
rect 547 -1761 577 -1721
rect 740 -1761 770 -1721
rect 900 -1761 930 -1721
rect 1100 -1761 1130 -1721
rect 1310 -1731 1330 -1691
rect 1370 -1731 1390 -1691
rect 387 -1781 427 -1761
rect 387 -1821 393 -1781
rect 423 -1821 427 -1781
rect 387 -1845 427 -1821
rect 467 -1781 507 -1761
rect 467 -1821 470 -1781
rect 500 -1821 507 -1781
rect 467 -1845 507 -1821
rect 547 -1781 587 -1761
rect 547 -1821 553 -1781
rect 583 -1821 587 -1781
rect 547 -1845 587 -1821
rect 627 -1781 667 -1761
rect 627 -1821 630 -1781
rect 660 -1821 667 -1781
rect 627 -1845 667 -1821
rect 740 -1781 780 -1761
rect 740 -1821 745 -1781
rect 776 -1821 780 -1781
rect 740 -1845 780 -1821
rect 818 -1781 858 -1761
rect 818 -1821 824 -1781
rect 854 -1821 858 -1781
rect 818 -1845 858 -1821
rect 900 -1781 940 -1761
rect 900 -1821 906 -1781
rect 936 -1821 940 -1781
rect 900 -1845 940 -1821
rect 980 -1781 1020 -1761
rect 980 -1821 985 -1781
rect 1015 -1821 1020 -1781
rect 980 -1845 1020 -1821
rect 1100 -1781 1140 -1761
rect 1100 -1821 1106 -1781
rect 1136 -1821 1140 -1781
rect 1100 -1845 1140 -1821
rect 1180 -1781 1220 -1761
rect 1180 -1821 1183 -1781
rect 1213 -1821 1220 -1781
rect 1180 -1845 1220 -1821
rect 12 -1991 52 -1981
rect -30 -2011 22 -1991
rect 42 -2011 52 -1991
rect -30 -2021 52 -2011
rect 77 -2121 107 -1845
rect 228 -1942 258 -1845
rect 277 -1891 317 -1881
rect 277 -1911 287 -1891
rect 307 -1911 317 -1891
rect 277 -1921 317 -1911
rect 407 -1942 447 -1932
rect 228 -1962 417 -1942
rect 437 -1962 447 -1942
rect 228 -1972 447 -1962
rect 249 -2078 292 -2071
rect 249 -2105 258 -2078
rect 284 -2105 292 -2078
rect 249 -2114 292 -2105
rect 77 -2131 212 -2121
rect 77 -2151 182 -2131
rect 202 -2151 212 -2131
rect 77 -2269 107 -2151
rect 172 -2161 212 -2151
rect 312 -2227 342 -1972
rect -13 -2279 27 -2269
rect -13 -2303 -5 -2279
rect 19 -2303 27 -2279
rect -13 -2311 27 -2303
rect 67 -2279 107 -2269
rect 67 -2303 75 -2279
rect 99 -2303 107 -2279
rect 67 -2311 107 -2303
rect 147 -2235 187 -2227
rect 147 -2303 155 -2235
rect 179 -2303 187 -2235
rect 147 -2311 187 -2303
rect 302 -2235 342 -2227
rect 302 -2303 311 -2235
rect 335 -2303 342 -2235
rect 477 -1991 507 -1845
rect 637 -1941 667 -1845
rect 823 -1881 853 -1845
rect 990 -1881 1020 -1845
rect 820 -1891 1020 -1881
rect 820 -1911 830 -1891
rect 850 -1911 1020 -1891
rect 820 -1921 860 -1911
rect 637 -1951 800 -1941
rect 637 -1971 770 -1951
rect 790 -1971 800 -1951
rect 477 -2001 607 -1991
rect 477 -2021 577 -2001
rect 597 -2021 607 -2001
rect 477 -2269 507 -2021
rect 567 -2031 607 -2021
rect 637 -2269 667 -1971
rect 760 -1981 800 -1971
rect 842 -2028 885 -2021
rect 842 -2055 851 -2028
rect 877 -2055 885 -2028
rect 842 -2064 885 -2055
rect 904 -2081 934 -1911
rect 1190 -1931 1220 -1845
rect 1310 -1771 1390 -1731
rect 1310 -1811 1330 -1771
rect 1370 -1811 1390 -1771
rect 1310 -1851 1390 -1811
rect 1310 -1891 1330 -1851
rect 1370 -1891 1390 -1851
rect 1310 -1931 1390 -1891
rect 1190 -1961 1260 -1931
rect 955 -1988 998 -1981
rect 955 -2015 964 -1988
rect 990 -2015 998 -1988
rect 955 -2024 998 -2015
rect 730 -2088 934 -2081
rect 730 -2114 737 -2088
rect 763 -2111 934 -2088
rect 763 -2114 770 -2111
rect 730 -2121 770 -2114
rect 904 -2121 934 -2111
rect 1125 -2121 1165 -2111
rect 904 -2141 1135 -2121
rect 1155 -2141 1165 -2121
rect 904 -2151 1165 -2141
rect 980 -2185 1010 -2151
rect 302 -2311 342 -2303
rect 387 -2279 427 -2269
rect 387 -2303 395 -2279
rect 419 -2303 427 -2279
rect 387 -2311 427 -2303
rect 467 -2279 507 -2269
rect 467 -2303 475 -2279
rect 499 -2303 507 -2279
rect 467 -2311 507 -2303
rect 547 -2279 587 -2269
rect 547 -2303 555 -2279
rect 579 -2303 587 -2279
rect 547 -2311 587 -2303
rect 627 -2279 667 -2269
rect 627 -2303 635 -2279
rect 659 -2303 667 -2279
rect 627 -2311 667 -2303
rect 740 -2221 780 -2185
rect 740 -2289 748 -2221
rect 772 -2289 780 -2221
rect 740 -2311 780 -2289
rect 980 -2212 1020 -2185
rect 980 -2280 988 -2212
rect 1012 -2280 1020 -2212
rect 1190 -2269 1220 -1961
rect 980 -2311 1020 -2280
rect 1100 -2279 1140 -2269
rect 1100 -2303 1108 -2279
rect 1132 -2303 1140 -2279
rect 1100 -2311 1140 -2303
rect 1180 -2279 1220 -2269
rect 1180 -2303 1188 -2279
rect 1212 -2303 1220 -2279
rect 1180 -2311 1220 -2303
rect 1310 -1971 1330 -1931
rect 1370 -1971 1390 -1931
rect 1310 -2011 1390 -1971
rect 1310 -2051 1330 -2011
rect 1370 -2051 1390 -2011
rect 1310 -2091 1390 -2051
rect 1310 -2131 1330 -2091
rect 1370 -2131 1390 -2091
rect 1310 -2261 1390 -2131
rect 1310 -2301 1330 -2261
rect 1370 -2301 1390 -2261
rect -13 -2350 17 -2311
rect 147 -2350 177 -2311
rect 387 -2350 417 -2311
rect 547 -2350 577 -2311
rect 740 -2350 770 -2311
rect 1100 -2350 1130 -2311
rect 1310 -2350 1390 -2301
rect -70 -2370 1390 -2350
rect -70 -2410 -40 -2370
rect 0 -2410 40 -2370
rect 80 -2410 120 -2370
rect 160 -2410 200 -2370
rect 240 -2410 280 -2370
rect 320 -2410 360 -2370
rect 400 -2410 440 -2370
rect 480 -2410 520 -2370
rect 560 -2410 600 -2370
rect 640 -2410 680 -2370
rect 720 -2410 760 -2370
rect 800 -2410 840 -2370
rect 880 -2410 920 -2370
rect 960 -2410 1000 -2370
rect 1040 -2410 1080 -2370
rect 1120 -2410 1160 -2370
rect 1200 -2410 1240 -2370
rect 1280 -2410 1320 -2370
rect 1360 -2410 1390 -2370
rect -70 -2430 1390 -2410
<< viali >>
rect 261 297 287 324
rect 290 110 310 130
rect 707 307 733 333
rect 821 247 847 274
rect 934 207 960 234
rect 800 110 820 130
rect 232 0 262 40
rect 375 -360 405 -320
rect 1056 -359 1086 -319
rect 320 -550 346 -524
rect 584 -600 606 -580
rect 1000 -550 1026 -524
rect 844 -600 866 -580
rect 920 -670 946 -644
rect 1080 -670 1106 -644
rect 1137 -897 1163 -776
rect 458 -1172 484 -1104
rect 1136 -1138 1162 -1112
rect 320 -1267 346 -1241
rect 320 -1377 346 -1351
rect 584 -1401 606 -1381
rect 1051 -1453 1077 -1427
rect 375 -1581 405 -1541
rect 229 -1821 259 -1781
rect 287 -1911 307 -1891
rect 258 -2105 284 -2078
rect 830 -1911 850 -1891
rect 851 -2055 877 -2028
rect 964 -2015 990 -1988
rect 737 -2114 763 -2088
<< metal1 >>
rect 700 333 740 340
rect 252 324 295 333
rect 252 297 261 324
rect 287 297 295 324
rect 700 307 707 333
rect 733 307 740 333
rect 700 300 740 307
rect 252 290 295 297
rect 812 274 855 283
rect 812 247 821 274
rect 847 247 855 274
rect 812 240 855 247
rect 925 234 968 243
rect 925 207 934 234
rect 960 207 968 234
rect 925 200 968 207
rect 280 130 320 140
rect 790 130 830 140
rect 280 110 290 130
rect 310 110 800 130
rect 820 110 830 130
rect 280 100 830 110
rect 227 40 267 64
rect 227 0 232 40
rect 262 0 267 40
rect 227 -20 267 0
rect 370 -320 410 -300
rect 370 -360 375 -320
rect 405 -360 410 -320
rect 370 -384 410 -360
rect 1050 -319 1090 -300
rect 1050 -359 1056 -319
rect 1086 -359 1090 -319
rect 1050 -384 1090 -359
rect 310 -524 355 -510
rect 310 -550 320 -524
rect 346 -550 355 -524
rect 310 -560 355 -550
rect 990 -524 1035 -510
rect 990 -550 1000 -524
rect 1026 -550 1035 -524
rect 990 -560 1035 -550
rect 575 -580 615 -570
rect 835 -580 875 -570
rect 575 -600 584 -580
rect 606 -600 844 -580
rect 866 -600 875 -580
rect 575 -610 875 -600
rect 910 -644 955 -630
rect 910 -670 920 -644
rect 946 -670 955 -644
rect 910 -680 955 -670
rect 1070 -644 1115 -630
rect 1070 -670 1080 -644
rect 1106 -670 1115 -644
rect 1070 -680 1115 -670
rect 1129 -776 1171 -748
rect 1129 -897 1137 -776
rect 1163 -897 1171 -776
rect 1129 -917 1171 -897
rect 450 -1104 492 -1094
rect 450 -1172 458 -1104
rect 484 -1172 492 -1104
rect 1128 -1112 1170 -1105
rect 1128 -1138 1136 -1112
rect 1162 -1138 1170 -1112
rect 1128 -1146 1170 -1138
rect 450 -1180 492 -1172
rect 310 -1241 355 -1231
rect 310 -1267 320 -1241
rect 346 -1267 355 -1241
rect 310 -1281 355 -1267
rect 310 -1351 355 -1341
rect 310 -1377 320 -1351
rect 346 -1377 355 -1351
rect 310 -1391 355 -1377
rect 575 -1381 615 -1371
rect 575 -1401 584 -1381
rect 606 -1401 615 -1381
rect 575 -1411 615 -1401
rect 1043 -1427 1085 -1420
rect 1043 -1453 1051 -1427
rect 1077 -1453 1085 -1427
rect 1043 -1461 1085 -1453
rect 370 -1541 410 -1517
rect 370 -1581 375 -1541
rect 405 -1581 410 -1541
rect 370 -1601 410 -1581
rect 224 -1781 264 -1761
rect 224 -1821 229 -1781
rect 259 -1821 264 -1781
rect 224 -1845 264 -1821
rect 277 -1891 860 -1881
rect 277 -1911 287 -1891
rect 307 -1911 830 -1891
rect 850 -1911 860 -1891
rect 277 -1921 317 -1911
rect 820 -1921 860 -1911
rect 955 -1988 998 -1981
rect 955 -2015 964 -1988
rect 990 -2015 998 -1988
rect 842 -2028 885 -2021
rect 955 -2024 998 -2015
rect 842 -2055 851 -2028
rect 877 -2055 885 -2028
rect 842 -2064 885 -2055
rect 249 -2078 292 -2071
rect 249 -2105 258 -2078
rect 284 -2105 292 -2078
rect 249 -2114 292 -2105
rect 730 -2088 770 -2081
rect 730 -2114 737 -2088
rect 763 -2114 770 -2088
rect 730 -2121 770 -2114
<< via1 >>
rect 261 297 287 324
rect 707 307 733 333
rect 821 247 847 274
rect 934 207 960 234
rect 232 0 262 40
rect 375 -360 405 -320
rect 1056 -359 1086 -319
rect 320 -550 346 -524
rect 1000 -550 1026 -524
rect 920 -670 946 -644
rect 1080 -670 1106 -644
rect 1137 -897 1163 -776
rect 458 -1172 484 -1104
rect 1136 -1138 1162 -1112
rect 320 -1267 346 -1241
rect 320 -1377 346 -1351
rect 1051 -1453 1077 -1427
rect 375 -1581 405 -1541
rect 229 -1821 259 -1781
rect 964 -2015 990 -1988
rect 851 -2055 877 -2028
rect 258 -2105 284 -2078
rect 737 -2114 763 -2088
<< metal2 >>
rect 700 333 740 340
rect 252 324 707 333
rect 252 297 261 324
rect 287 307 707 324
rect 733 307 740 333
rect 287 303 740 307
rect 287 297 295 303
rect 700 300 740 303
rect 252 290 295 297
rect 812 274 855 283
rect 812 270 821 274
rect 690 247 821 270
rect 847 247 855 274
rect 690 240 855 247
rect 227 40 267 64
rect 227 0 232 40
rect 262 0 267 40
rect 227 -20 267 0
rect 230 -520 260 -20
rect 690 -140 720 240
rect 925 234 968 243
rect 925 207 934 234
rect 960 230 968 234
rect 960 207 1040 230
rect 925 200 1040 207
rect 375 -170 720 -140
rect 1010 -140 1040 200
rect 1010 -170 1080 -140
rect 375 -300 405 -170
rect 1050 -300 1080 -170
rect 370 -320 410 -300
rect 370 -360 375 -320
rect 405 -360 410 -320
rect 370 -384 410 -360
rect 1050 -319 1090 -300
rect 1050 -359 1056 -319
rect 1086 -359 1090 -319
rect 1050 -384 1090 -359
rect 310 -520 355 -510
rect 990 -520 1035 -510
rect 230 -524 1035 -520
rect 230 -550 320 -524
rect 346 -550 1000 -524
rect 1026 -550 1035 -524
rect 310 -560 355 -550
rect 990 -560 1035 -550
rect 910 -644 955 -630
rect 910 -650 920 -644
rect 770 -670 920 -650
rect 946 -670 955 -644
rect 770 -680 955 -670
rect 1070 -644 1240 -630
rect 1070 -670 1080 -644
rect 1106 -660 1240 -644
rect 1106 -670 1115 -660
rect 1070 -680 1115 -670
rect 770 -986 800 -680
rect 462 -1016 800 -986
rect 1129 -776 1171 -748
rect 1129 -897 1137 -776
rect 1163 -897 1171 -776
rect 1129 -917 1171 -897
rect 462 -1094 492 -1016
rect 450 -1104 492 -1094
rect 450 -1172 458 -1104
rect 484 -1172 492 -1104
rect 1129 -1105 1159 -917
rect 1128 -1112 1170 -1105
rect 1128 -1138 1136 -1112
rect 1162 -1138 1170 -1112
rect 1128 -1146 1170 -1138
rect 450 -1180 492 -1172
rect 310 -1241 355 -1231
rect 310 -1267 320 -1241
rect 346 -1251 355 -1241
rect 1210 -1251 1240 -660
rect 346 -1267 1240 -1251
rect 310 -1281 1240 -1267
rect 310 -1351 355 -1341
rect 227 -1377 320 -1351
rect 346 -1377 355 -1351
rect 227 -1381 355 -1377
rect 227 -1761 257 -1381
rect 310 -1391 355 -1381
rect 1043 -1427 1085 -1420
rect 1043 -1453 1051 -1427
rect 1077 -1453 1085 -1427
rect 1043 -1461 1085 -1453
rect 370 -1541 410 -1517
rect 370 -1581 375 -1541
rect 405 -1581 410 -1541
rect 370 -1601 410 -1581
rect 375 -1671 405 -1601
rect 375 -1701 720 -1671
rect 224 -1781 264 -1761
rect 224 -1821 229 -1781
rect 259 -1821 264 -1781
rect 224 -1845 264 -1821
rect 690 -2021 720 -1701
rect 1050 -1981 1080 -1461
rect 955 -1988 1080 -1981
rect 955 -2015 964 -1988
rect 990 -2011 1080 -1988
rect 990 -2015 998 -2011
rect 690 -2028 885 -2021
rect 955 -2024 998 -2015
rect 690 -2051 851 -2028
rect 842 -2055 851 -2051
rect 877 -2055 885 -2028
rect 842 -2064 885 -2055
rect 249 -2078 292 -2071
rect 249 -2105 258 -2078
rect 284 -2084 292 -2078
rect 730 -2084 770 -2081
rect 284 -2088 770 -2084
rect 284 -2105 737 -2088
rect 249 -2114 737 -2105
rect 763 -2114 770 -2088
rect 730 -2121 770 -2114
<< labels >>
rlabel locali 1230 -1951 1250 -1941 1 dn
rlabel locali -20 -2011 0 -2001 1 fvco_8
rlabel locali 1340 -996 1360 -986 1 gnd!
rlabel locali -100 -906 -80 -886 1 vdd
rlabel locali 1200 160 1220 170 1 up
rlabel locali -20 210 0 220 1 fin
<< end >>
