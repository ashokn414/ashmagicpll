magic
tech sky130A
timestamp 1604917003
<< nwell >>
rect -87 -20 121 139
<< nmos >>
rect 0 -117 40 -75
<< pmos >>
rect 0 0 40 42
<< ndiff >>
rect -40 -84 0 -75
rect -40 -109 -35 -84
rect -15 -109 0 -84
rect -40 -117 0 -109
rect 40 -84 80 -75
rect 40 -109 55 -84
rect 75 -109 80 -84
rect 40 -117 80 -109
<< pdiff >>
rect -40 33 0 42
rect -40 8 -35 33
rect -15 8 0 33
rect -40 0 0 8
rect 40 33 80 42
rect 40 8 55 33
rect 75 8 80 33
rect 40 0 80 8
<< ndiffc >>
rect -35 -109 -15 -84
rect 55 -109 75 -84
<< pdiffc >>
rect -35 8 -15 33
rect 55 8 75 33
<< psubdiff >>
rect -58 -191 -15 -170
rect 6 -191 31 -170
rect 52 -191 86 -170
<< nsubdiff >>
rect -59 99 -23 120
rect -2 99 22 120
rect 43 99 86 120
<< psubdiffcont >>
rect -15 -191 6 -170
rect 31 -191 52 -170
<< nsubdiffcont >>
rect -23 99 -2 120
rect 22 99 43 120
<< poly >>
rect 0 42 40 67
rect 0 -25 40 0
rect -35 -31 40 -25
rect -35 -49 -25 -31
rect -8 -49 40 -31
rect -35 -58 40 -49
rect 0 -75 40 -58
rect 0 -137 40 -117
<< polycont >>
rect -25 -49 -8 -31
<< locali >>
rect -70 120 102 125
rect -70 99 -54 120
rect -33 99 22 120
rect 43 99 57 120
rect 78 99 102 120
rect -70 95 102 99
rect -40 33 -15 95
rect -40 8 -35 33
rect -40 0 -15 8
rect 55 33 80 42
rect 75 8 80 33
rect -35 -31 0 -25
rect -35 -49 -25 -31
rect -8 -49 0 -31
rect -35 -58 0 -49
rect -40 -84 -15 -75
rect -40 -109 -35 -84
rect -40 -162 -15 -109
rect 55 -84 80 8
rect 75 -109 80 -84
rect 55 -117 80 -109
rect -70 -170 100 -162
rect -70 -191 -51 -170
rect -30 -191 -15 -170
rect 6 -191 31 -170
rect 52 -191 63 -170
rect 84 -191 100 -170
rect -70 -197 100 -191
<< viali >>
rect -54 99 -33 120
rect 57 99 78 120
rect -51 -191 -30 -170
rect 63 -191 84 -170
<< metal1 >>
rect -83 120 115 131
rect -83 99 -54 120
rect -33 99 57 120
rect 78 99 115 120
rect -83 88 115 99
rect -83 -170 115 -157
rect -83 -191 -51 -170
rect -30 -191 63 -170
rect 84 -191 115 -170
rect -83 -201 115 -191
<< labels >>
flabel locali s -25 -49 -8 -31 0 FreeSans 120 0 0 0 A
port 1 nsew
flabel locali s 55 -50 80 -30 0 FreeSans 120 0 0 0 Y
port 3 nsew
flabel metal1 s -10 98 56 114 0 FreeSans 120 0 0 0 VPWR
port 5 nsew
flabel metal1 s -13 -182 44 -166 0 FreeSans 120 0 0 0 VGND
port 6 nsew
<< end >>
